
module remap ( m1, m2 );
  input [27:0] m1;
  output [26:0] m2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n121, n122, n123,
         n124, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n175, n176, n177, n179, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n199, n200, n201, n202, n203, n204, n205,
         n206, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n223, n224, n225, n226, n227, n228, n230,
         n231, n232, n233, n234, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1170, n1171, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042;

  AN2BSVTX2 U3 ( .A(n1308), .B(n1563), .Z(n1313) );
  IVSVTX0H U4 ( .A(n1945), .Z(n1968) );
  AO2SVTX1 U5 ( .A(n1718), .B(n1901), .C(n165), .D(n772), .Z(n1902) );
  AO6SVTX1 U6 ( .A(n543), .B(n1470), .C(n1469), .Z(n1471) );
  ND2SVTX2 U7 ( .A(n402), .B(n697), .Z(n155) );
  NR2SVTX2 U8 ( .A(n1975), .B(n197), .Z(n1976) );
  NR2SVTX1 U9 ( .A(n444), .B(n1652), .Z(n1476) );
  ENSVTX1 U10 ( .A(n1740), .B(n1739), .Z(n1794) );
  AO2SVTX2 U11 ( .A(n1818), .B(n1488), .C(n1817), .D(n1718), .Z(n1834) );
  AO6SVTX1 U12 ( .A(n102), .B(n742), .C(n1316), .Z(n1317) );
  NR2ASVTX1 U13 ( .A(n1579), .B(n1578), .Z(n1587) );
  ND2ASVTX6 U14 ( .A(n92), .B(n1573), .Z(n1979) );
  ND3SVTX2 U15 ( .A(n1375), .B(n1374), .C(n1373), .Z(n1376) );
  NR2ASVTX1 U16 ( .A(n1796), .B(n1795), .Z(n1801) );
  OR2SVTX1 U17 ( .A(n1192), .B(n1191), .Z(n697) );
  NR2ASVTX1 U18 ( .A(n45), .B(n1737), .Z(n1740) );
  IVSVTX0H U19 ( .A(n334), .Z(n1611) );
  BFSVTX2 U20 ( .A(n2029), .Z(n128) );
  IVSVTX2 U21 ( .A(n22), .Z(n1507) );
  EOSVTX0H U22 ( .A(n1778), .B(n1777), .Z(n1791) );
  CTBUFSVTX4 U23 ( .A(n398), .Z(n212) );
  IVSVTX0H U24 ( .A(n1994), .Z(n1798) );
  IVSVTX2 U25 ( .A(n1539), .Z(n202) );
  IVSVTX0H U26 ( .A(n143), .Z(n505) );
  CTIVSVTX2 U27 ( .A(n1973), .Z(n1975) );
  AN2BSVTX2 U28 ( .A(n1963), .B(n2029), .Z(n1964) );
  AO6SVTX1 U29 ( .A(n1320), .B(n1986), .C(n1985), .Z(n1987) );
  NR2ASVTX1 U30 ( .A(n1443), .B(n7), .Z(n1702) );
  IVSVTX2 U31 ( .A(n225), .Z(n1322) );
  CTAN2BSVTX4 U32 ( .A(n1540), .B(n1549), .Z(n1538) );
  B_ND2SVTX1 U33 ( .A(n806), .B(n372), .Z(n1373) );
  OR2BSVTX4 U34 ( .A(n690), .B(n1646), .Z(n1971) );
  NR2ASVTX1 U35 ( .A(n1607), .B(n901), .Z(n334) );
  BFSVTX0H U36 ( .A(n1441), .Z(n7) );
  IVSVTX0H U37 ( .A(n1909), .Z(n1911) );
  CTIVSVTX2 U38 ( .A(n1552), .Z(n184) );
  IVSVTX0H U39 ( .A(n1634), .Z(n1636) );
  IVSVTX0H U40 ( .A(n1694), .Z(n1897) );
  IVSVTX0H U41 ( .A(n1873), .Z(n1874) );
  IVSVTX0H U42 ( .A(n1688), .Z(n1877) );
  BFSVTX0H U43 ( .A(n1693), .Z(n138) );
  IVSVTX0H U44 ( .A(n1805), .Z(n1806) );
  IVSVTX0H U45 ( .A(n753), .Z(n1840) );
  IVSVTX0H U46 ( .A(n1719), .Z(n1720) );
  IVSVTX2 U47 ( .A(n1652), .Z(n420) );
  AO6SVTX1 U48 ( .A(n1656), .B(n276), .C(n1727), .Z(n1728) );
  BFSVTX0H U49 ( .A(n1608), .Z(n151) );
  IVSVTX0H U50 ( .A(n1658), .Z(n1723) );
  IVSVTX0H U51 ( .A(n682), .Z(n1714) );
  IVSVTX0H U52 ( .A(n1401), .Z(n1402) );
  IVSVTX0H U53 ( .A(n1668), .Z(n1708) );
  CTBUFSVTX2 U54 ( .A(n568), .Z(n169) );
  IVSVTX0H U55 ( .A(n9), .Z(n1379) );
  IVSVTX0H U56 ( .A(n1360), .Z(n1319) );
  IVSVTX0H U57 ( .A(n1600), .Z(n1601) );
  IVSVTX0H U58 ( .A(n722), .Z(n852) );
  IVSVTX0H U59 ( .A(n1984), .Z(n1985) );
  IVSVTX0H U60 ( .A(n1395), .Z(n506) );
  IVSVTX0H U61 ( .A(n1614), .Z(n1616) );
  IVSVTX0H U62 ( .A(n589), .Z(n762) );
  NR2SVTX8 U63 ( .A(n1795), .B(n1799), .Z(n1915) );
  IVSVTX0H U64 ( .A(n156), .Z(n1451) );
  IVSVTX0H U65 ( .A(n164), .Z(n1458) );
  IVSVTX0H U66 ( .A(n1983), .Z(n1986) );
  IVSVTX0H U67 ( .A(n1419), .Z(n725) );
  AN2SVTX0H U68 ( .A(n140), .B(n433), .Z(n685) );
  NR2SVTX6 U69 ( .A(n1563), .B(n1653), .Z(n396) );
  IVSVTX0H U70 ( .A(n154), .Z(n1814) );
  IVSVTX0H U71 ( .A(n981), .Z(n965) );
  IVSVTX0H U72 ( .A(n1825), .Z(n1406) );
  IVSVTX2 U73 ( .A(n567), .Z(n1652) );
  IVSVTX0H U74 ( .A(n1912), .Z(n1913) );
  IVSVTX0H U75 ( .A(n1582), .Z(n1583) );
  BFSVTX0H U76 ( .A(n1773), .Z(n164) );
  BFSVTX0H U77 ( .A(n1759), .Z(n24) );
  BFSVTX0H U78 ( .A(n1744), .Z(n156) );
  BFSVTX0H U79 ( .A(n723), .Z(n154) );
  IVSVTX0H U80 ( .A(n1918), .Z(n1919) );
  IVSVTX4 U81 ( .A(n402), .Z(n92) );
  IVSVTX4 U82 ( .A(n1553), .Z(n1562) );
  NR2SVTX4 U83 ( .A(n1653), .B(n1563), .Z(n553) );
  IVSVTX0H U84 ( .A(n1365), .Z(n1366) );
  IVSVTX0H U85 ( .A(n1326), .Z(n1920) );
  BFSVTX0H U86 ( .A(n2034), .Z(n9) );
  IVSVTX0H U87 ( .A(n2032), .Z(n2035) );
  IVSVTX2 U88 ( .A(n244), .Z(n34) );
  IVSVTX0H U89 ( .A(n2004), .Z(n2006) );
  CTIVSVTX2 U90 ( .A(n1993), .Z(n693) );
  IVSVTX0H U91 ( .A(n1463), .Z(n1466) );
  IVSVTX0H U92 ( .A(n2014), .Z(n2022) );
  CTBUFSVTX2 U93 ( .A(n1756), .Z(n23) );
  IVSVTX0H U94 ( .A(n1664), .Z(n1435) );
  IVSVTX0H U95 ( .A(n1663), .Z(n1436) );
  BFSVTX0H U96 ( .A(n1726), .Z(n47) );
  AO7SVTX6 U97 ( .A(n939), .B(n358), .C(n37), .Z(n1549) );
  IVSVTX2 U98 ( .A(n26), .Z(n624) );
  NR2ASVTX4 U99 ( .A(n718), .B(n1094), .Z(n389) );
  ND2ASVTX4 U100 ( .A(n1146), .B(n1193), .Z(n1973) );
  IVSVTX0H U101 ( .A(n1513), .Z(n1514) );
  CTIVSVTX4 U102 ( .A(n1645), .Z(n1646) );
  IVSVTX0H U103 ( .A(n333), .Z(n2018) );
  CTIVSVTX2 U104 ( .A(n1284), .Z(n658) );
  ND2SVTX2 U105 ( .A(n67), .B(n1488), .Z(n39) );
  ND3SVTX6 U106 ( .A(n1118), .B(n69), .C(n490), .Z(n1083) );
  IVSVTX0H U107 ( .A(n972), .Z(n1438) );
  ND3ABSVTX2 U108 ( .A(n1463), .B(n1327), .C(n1462), .Z(n1328) );
  BFSVTX2 U109 ( .A(n938), .Z(n37) );
  CTIVSVTX2 U110 ( .A(n994), .Z(n995) );
  ND2ASVTX6 U111 ( .A(n1597), .B(n451), .Z(n415) );
  IVSVTX2 U112 ( .A(n295), .Z(n126) );
  CTIVSVTX2 U113 ( .A(n1194), .Z(n1146) );
  IVSVTX0H U114 ( .A(n993), .Z(n996) );
  IVSVTX2 U115 ( .A(n1095), .Z(n590) );
  ND2SVTX2 U116 ( .A(n1141), .B(n1488), .Z(n417) );
  NR2SVTX6 U117 ( .A(n241), .B(n1483), .Z(n240) );
  OR2SVTX1 U118 ( .A(n1245), .B(n1145), .Z(n292) );
  AO6SVTX6 U119 ( .A(n1063), .B(n543), .C(n176), .Z(n1064) );
  ND2SVTX2 U120 ( .A(n168), .B(n728), .Z(n472) );
  CTBUFSVTX6 U121 ( .A(n281), .Z(n718) );
  ND2ASVTX6 U122 ( .A(n1597), .B(n301), .Z(n300) );
  IVSVTX10 U123 ( .A(n1488), .Z(n81) );
  IVSVTX0H U124 ( .A(n1144), .Z(n1245) );
  NR2SVTX2 U125 ( .A(n669), .B(n13), .Z(n836) );
  NR2SVTX4 U126 ( .A(n487), .B(n281), .Z(n295) );
  NR2ASVTX2 U127 ( .A(n1087), .B(n82), .Z(n1086) );
  ND3SVTX4 U128 ( .A(n336), .B(n1164), .C(n265), .Z(n54) );
  AN2SVTX2 U129 ( .A(n674), .B(n1119), .Z(n766) );
  BFSVTX0H U130 ( .A(m1[25]), .Z(n129) );
  ND2ASVTX6 U131 ( .A(n1175), .B(n806), .Z(n620) );
  IVSVTX2 U132 ( .A(n1084), .Z(n137) );
  IVSVTX0H U133 ( .A(n119), .Z(n211) );
  IVSVTX2 U134 ( .A(n1240), .Z(n13) );
  ND2SVTX2 U135 ( .A(n715), .B(n1164), .Z(n621) );
  IVSVTX6 U136 ( .A(n1597), .Z(n543) );
  ND2SVTX2 U137 ( .A(n872), .B(n362), .Z(n878) );
  ND3SVTX6 U138 ( .A(n434), .B(n1087), .C(n466), .Z(n1062) );
  AO6SVTX6 U139 ( .A(n74), .B(n1116), .C(n1115), .Z(n1117) );
  ND3SVTX4 U140 ( .A(n96), .B(n631), .C(n987), .Z(n359) );
  ND3SVTX4 U141 ( .A(n876), .B(n873), .C(n1008), .Z(n879) );
  NR3ABSVTX4 U142 ( .A(n106), .B(n717), .C(n1280), .Z(n1490) );
  ND3ABSVTX2 U143 ( .A(n730), .B(n1295), .C(n1286), .Z(n1285) );
  NR2SVTX2 U144 ( .A(n717), .B(n674), .Z(n48) );
  AN2SVTX1 U145 ( .A(n1187), .B(n204), .Z(n1188) );
  NR2SVTX2 U146 ( .A(n728), .B(n135), .Z(n481) );
  IVSVTX2 U147 ( .A(n1119), .Z(n710) );
  IVSVTX2 U148 ( .A(n1009), .Z(n602) );
  BFSVTX8 U149 ( .A(n1275), .Z(n467) );
  ND2ASVTX6 U150 ( .A(n660), .B(n1482), .Z(n1087) );
  NR2SVTX2 U151 ( .A(n804), .B(n492), .Z(n988) );
  IVSVTX0H U152 ( .A(n1127), .Z(n113) );
  BFSVTX0H U153 ( .A(n1080), .Z(n57) );
  CTIVSVTX2 U154 ( .A(n1012), .Z(n1559) );
  IVSVTX0H U155 ( .A(n1031), .Z(n1032) );
  IVSVTX0H U156 ( .A(n1241), .Z(n135) );
  BFSVTX6 U157 ( .A(n1259), .Z(n1320) );
  IVSVTX0H U158 ( .A(n1129), .Z(n1162) );
  ND3ASVTX4 U159 ( .A(n789), .B(n366), .C(n365), .Z(n1499) );
  BFSVTX4 U160 ( .A(n1111), .Z(n8) );
  IVSVTX2 U161 ( .A(n215), .Z(n790) );
  CTIVSVTX2 U162 ( .A(n1502), .Z(n717) );
  NR2ASVTX4 U163 ( .A(n36), .B(n1517), .Z(n1504) );
  ND2SVTX2 U164 ( .A(n545), .B(n78), .Z(n936) );
  IVSVTX8 U165 ( .A(n321), .Z(n306) );
  ND2SVTX2 U166 ( .A(n1484), .B(n876), .Z(n874) );
  IVSVTX6 U167 ( .A(n675), .Z(n299) );
  ND2ASVTX6 U168 ( .A(n227), .B(n230), .Z(n434) );
  BFSVTX0H U169 ( .A(n915), .Z(n215) );
  CTIVSVTX2 U170 ( .A(n1494), .Z(n1295) );
  IVSVTX6 U171 ( .A(n345), .Z(n96) );
  IVSVTX2 U172 ( .A(n1048), .Z(n1049) );
  IVSVTX0H U173 ( .A(n1052), .Z(n1053) );
  ND2SVTX6 U174 ( .A(n937), .B(n1167), .Z(n728) );
  IVSVTX2 U175 ( .A(n1182), .Z(n1075) );
  NR2ASVTX4 U176 ( .A(n1287), .B(n1492), .Z(n1293) );
  IVSVTX0H U177 ( .A(n1199), .Z(n1200) );
  OR2SVTX2 U178 ( .A(n1197), .B(n837), .Z(n1012) );
  IVSVTX0H U179 ( .A(n1104), .Z(n1035) );
  ND2ASVTX6 U180 ( .A(n1011), .B(n1009), .Z(n403) );
  IVSVTX0H U181 ( .A(n1502), .Z(n36) );
  IVSVTX0H U182 ( .A(n757), .Z(n243) );
  B_ND2SVTX2 U183 ( .A(n1070), .B(n1069), .Z(n1076) );
  IVSVTX2 U184 ( .A(n928), .Z(n441) );
  ND2SVTX2 U185 ( .A(n1072), .B(n1071), .Z(n1143) );
  IVSVTX4 U186 ( .A(n517), .Z(n1074) );
  IVSVTX0H U187 ( .A(n551), .Z(n208) );
  ND2SVTX4 U188 ( .A(n937), .B(n1167), .Z(n1627) );
  IVSVTX4 U189 ( .A(n652), .Z(n634) );
  BFSVTX6 U190 ( .A(n1394), .Z(n563) );
  NR2SVTX2 U191 ( .A(n168), .B(n1529), .Z(n998) );
  IVSVTX2 U192 ( .A(n555), .Z(n1010) );
  AO7SVTX1 U193 ( .A(n569), .B(n1984), .C(n1982), .Z(n1211) );
  F_ND2ASVTX2 U194 ( .A(n177), .B(n796), .Z(n1069) );
  NR3SVTX6 U195 ( .A(n108), .B(n666), .C(n1264), .Z(n1136) );
  AO6SVTX4 U196 ( .A(n1991), .B(n56), .C(n1220), .Z(n1227) );
  ND4ABSVTX6 U197 ( .A(n449), .B(n1515), .C(n1242), .D(n1513), .Z(n210) );
  IVSVTX2 U198 ( .A(n1989), .Z(n1991) );
  CTIVSVTX2 U199 ( .A(n1045), .Z(n111) );
  IVSVTX2 U200 ( .A(n1100), .Z(n79) );
  ND2SVTX4 U201 ( .A(n1954), .B(n932), .Z(n410) );
  ND4ABSVTX6 U202 ( .A(n789), .B(n1171), .C(n847), .D(n261), .Z(n230) );
  IVSVTX2 U203 ( .A(n1981), .Z(n569) );
  IVSVTX4 U204 ( .A(n1228), .Z(n1993) );
  BFSVTX6 U205 ( .A(n767), .Z(n532) );
  CTIVSVTX2 U206 ( .A(n250), .Z(n1097) );
  AO3CDSVTX6 U207 ( .A(n1071), .B(n1072), .C(n87), .D(n75), .Z(n323) );
  AO7SVTX4 U208 ( .A(n1114), .B(n1022), .C(n1023), .Z(n370) );
  ND4SVTX6 U209 ( .A(n644), .B(n645), .C(n646), .D(n643), .Z(n1341) );
  AO7ABSVTX2 U210 ( .A(n103), .B(n549), .C(n1015), .Z(n547) );
  ND2SVTX2 U211 ( .A(n910), .B(n916), .Z(n1023) );
  F_IVSVTX1 U212 ( .A(m1[25]), .Z(n911) );
  ND2SVTX2 U213 ( .A(n916), .B(n119), .Z(n1046) );
  NR2SVTX4 U214 ( .A(n1219), .B(n1218), .Z(n1989) );
  CTIVSVTX2 U215 ( .A(n810), .Z(n1166) );
  IVSVTX2 U216 ( .A(n487), .Z(n789) );
  IVSVTX2 U217 ( .A(n799), .Z(n554) );
  IVSVTX2 U218 ( .A(n1578), .Z(n647) );
  B_ND2SVTX2 U219 ( .A(n1251), .B(n1249), .Z(n1203) );
  IVSVTX0H U220 ( .A(n890), .Z(n442) );
  NR3ABSVTX2 U221 ( .A(m1[27]), .B(n910), .C(n448), .Z(n447) );
  AO7SVTX2 U222 ( .A(n540), .B(n883), .C(n168), .Z(n885) );
  IVSVTX1 U223 ( .A(n1197), .Z(n14) );
  NR2SVTX6 U224 ( .A(n981), .B(n1442), .Z(n1441) );
  AN2BSVTX2 U225 ( .A(n669), .B(m1[24]), .Z(n783) );
  ND2ASVTX6 U226 ( .A(m1[16]), .B(n114), .Z(n1952) );
  EN3SVTX6 U227 ( .A(n869), .B(n572), .C(n904), .Z(n801) );
  IVSVTX6 U228 ( .A(n653), .Z(n561) );
  AN2SVTX6 U229 ( .A(n119), .B(n168), .Z(n1494) );
  CTIVSVTX2 U230 ( .A(n1036), .Z(n1105) );
  NR2ASVTX4 U231 ( .A(n918), .B(n88), .Z(n1264) );
  NR2SVTX4 U232 ( .A(n1252), .B(n1246), .Z(n906) );
  NR2SVTX6 U233 ( .A(n1433), .B(n1432), .Z(n967) );
  AO7SVTX6 U234 ( .A(n1386), .B(n1909), .C(n1910), .Z(n1342) );
  ND2SVTX4 U235 ( .A(n1769), .B(n541), .Z(n925) );
  ND2SVTX2 U236 ( .A(n1395), .B(n1391), .Z(n259) );
  IVSVTX2 U237 ( .A(n1554), .Z(n1518) );
  NR3SVTX2 U238 ( .A(n819), .B(n456), .C(n971), .Z(n691) );
  IVSVTX2 U239 ( .A(n1263), .Z(n1) );
  IVSVTX2 U240 ( .A(n250), .Z(n25) );
  IVSVTX10 U241 ( .A(n910), .Z(n119) );
  IVSVTX2 U242 ( .A(n511), .Z(n510) );
  ND2ASVTX6 U243 ( .A(m1[13]), .B(n277), .Z(n1337) );
  ND2ASVTX6 U244 ( .A(n114), .B(n916), .Z(n1133) );
  ND2ASVTX6 U245 ( .A(n53), .B(n805), .Z(n279) );
  NR2ASVTX4 U246 ( .A(n572), .B(n807), .Z(n1246) );
  B_ND2SVTX2 U247 ( .A(n933), .B(n76), .Z(n1036) );
  IVSVTX2 U248 ( .A(n851), .Z(n361) );
  ND2SVTX2 U249 ( .A(n920), .B(n80), .Z(n1810) );
  CTIVSVTX2 U250 ( .A(n1500), .Z(n1554) );
  CTIVSVTX2 U251 ( .A(n655), .Z(n337) );
  ND2ASVTX4 U252 ( .A(m1[11]), .B(n355), .Z(n1391) );
  NR2SVTX4 U253 ( .A(n511), .B(n108), .Z(n809) );
  IVSVTX2 U254 ( .A(n1416), .Z(n605) );
  ND2ASVTX4 U255 ( .A(n887), .B(n888), .Z(n882) );
  NR2SVTX2 U256 ( .A(n1609), .B(n90), .Z(n723) );
  NR2SVTX4 U257 ( .A(n1223), .B(n962), .Z(n1799) );
  NR2SVTX6 U258 ( .A(n1767), .B(n1773), .Z(n541) );
  F_ND3SVTX2 U259 ( .A(n890), .B(n910), .C(n1529), .Z(n1016) );
  IVSVTX2 U260 ( .A(n2002), .Z(n15) );
  NR2SVTX2 U261 ( .A(m1[27]), .B(m1[25]), .Z(n881) );
  CTBUFSVTX8 U262 ( .A(n1140), .Z(n133) );
  IVSVTX2 U263 ( .A(m1[27]), .Z(n890) );
  ND2ASVTX6 U264 ( .A(n895), .B(n696), .Z(n1876) );
  IVSVTX2 U265 ( .A(n1592), .Z(n209) );
  IVSVTX2 U266 ( .A(n195), .Z(n944) );
  B_ND2SVTX2 U267 ( .A(n355), .B(n704), .Z(n1931) );
  IVSVTX2 U268 ( .A(n480), .Z(n479) );
  CTBUFSVTX4 U269 ( .A(n784), .Z(n2) );
  B_ND2SVTX2 U270 ( .A(n807), .B(n957), .Z(n1151) );
  ND2SVTX2 U271 ( .A(n917), .B(n114), .Z(n1256) );
  IVSVTX2 U272 ( .A(n280), .Z(n53) );
  CTIVSVTX2 U273 ( .A(n430), .Z(n426) );
  AN2SVTX6 U274 ( .A(n777), .B(n735), .Z(n901) );
  ND2SVTX2 U275 ( .A(n140), .B(n1837), .Z(n1846) );
  ND2SVTX6 U276 ( .A(n408), .B(n497), .Z(n414) );
  ND2SVTX2 U277 ( .A(n896), .B(n894), .Z(n382) );
  NR2SVTX4 U278 ( .A(n1744), .B(n1741), .Z(n607) );
  NR3SVTX4 U279 ( .A(n1140), .B(n957), .C(n76), .Z(n424) );
  F_IVSVTX1 U280 ( .A(m1[25]), .Z(n356) );
  B_ND2SVTX2 U281 ( .A(n920), .B(n947), .Z(n1935) );
  ND2ASVTX6 U282 ( .A(n704), .B(n89), .Z(n849) );
  B_ND2SVTX2 U283 ( .A(n80), .B(n777), .Z(n1802) );
  ND2SVTX2 U284 ( .A(n920), .B(n28), .Z(n1361) );
  ND2SVTX2 U285 ( .A(n405), .B(n947), .Z(n949) );
  IVSVTX2 U286 ( .A(n950), .Z(n131) );
  IVSVTX6 U287 ( .A(n593), .Z(n19) );
  CTIVSVTX2 U288 ( .A(n274), .Z(n58) );
  BFSVTX8 U289 ( .A(n699), .Z(n140) );
  IVSVTX10 U290 ( .A(n429), .Z(n592) );
  CTBUFSVTX4 U291 ( .A(n1358), .Z(n21) );
  ND2SVTX4 U292 ( .A(n1323), .B(n1326), .Z(n2013) );
  IVSVTX2 U293 ( .A(n1150), .Z(n109) );
  ND2ASVTX6 U294 ( .A(n525), .B(n585), .Z(n1937) );
  CTBUFSVTX4 U295 ( .A(n1836), .Z(n203) );
  ND2ASVTX4 U296 ( .A(n80), .B(n704), .Z(n1803) );
  CTIVSVTX2 U297 ( .A(n1885), .Z(n858) );
  AN2SVTX4 U298 ( .A(n920), .B(m1[16]), .Z(n903) );
  NR2ASVTX4 U299 ( .A(n28), .B(n838), .Z(n570) );
  ND2SVTX4 U300 ( .A(n572), .B(n153), .Z(n478) );
  ND2SVTX4 U301 ( .A(n333), .B(n535), .Z(n824) );
  IVSVTX8 U302 ( .A(n619), .Z(n107) );
  IVSVTX4 U303 ( .A(n1712), .Z(n381) );
  ND4ABSVTX6 U304 ( .A(n405), .B(n408), .C(n317), .D(n10), .Z(n247) );
  AO7SVTX4 U305 ( .A(n1403), .B(n1824), .C(n1401), .Z(n815) );
  ND2SVTX2 U306 ( .A(m1[11]), .B(m1[13]), .Z(n1401) );
  ND2ASVTX6 U307 ( .A(n705), .B(n353), .Z(n1712) );
  IVSVTX6 U308 ( .A(n1140), .Z(n114) );
  IVSVTX2 U309 ( .A(n704), .Z(n335) );
  BFSVTX8 U310 ( .A(n918), .Z(n121) );
  CTIVSVTX2 U311 ( .A(n460), .Z(n459) );
  BFSVTX4 U312 ( .A(n473), .Z(n10) );
  IVSVTX10 U313 ( .A(n791), .Z(n915) );
  ND2SVTX2 U314 ( .A(m1[11]), .B(n706), .Z(n1615) );
  B_ND2SVTX2 U315 ( .A(n588), .B(n572), .Z(n1982) );
  ND2ASVTX6 U316 ( .A(n31), .B(n30), .Z(n1623) );
  ND2SVTX6 U317 ( .A(n963), .B(n897), .Z(n1607) );
  IVSVTX4 U318 ( .A(n353), .Z(n32) );
  ND3SVTX6 U319 ( .A(n162), .B(n507), .C(n526), .Z(n839) );
  B_ND2SVTX2 U320 ( .A(n500), .B(n735), .Z(n499) );
  ND2ASVTX6 U321 ( .A(m1[3]), .B(n950), .Z(n460) );
  IVSVTX8 U322 ( .A(n572), .Z(n566) );
  IVSVTX4 U323 ( .A(n526), .Z(n167) );
  IVSVTX8 U324 ( .A(n918), .Z(n957) );
  IVSVTX8 U325 ( .A(n588), .Z(n393) );
  IVSVTX6 U326 ( .A(n699), .Z(n456) );
  IVSVTX10 U327 ( .A(m1[14]), .Z(n355) );
  F_EOSVTX2 U328 ( .A(m1[1]), .B(m1[3]), .Z(n1837) );
  IVSVTX8 U329 ( .A(n777), .Z(n704) );
  NR2SVTX2 U330 ( .A(n1836), .B(n391), .Z(n1870) );
  IVSVTX4 U331 ( .A(n527), .Z(n384) );
  IVSVTX4 U332 ( .A(n716), .Z(n317) );
  IVSVTX8 U333 ( .A(n473), .Z(n116) );
  BFSVTX6 U334 ( .A(m1[6]), .Z(n408) );
  IVSVTX4 U335 ( .A(n535), .Z(n817) );
  ND2SVTX4 U336 ( .A(n274), .B(n950), .Z(n1323) );
  IVSVTX4 U337 ( .A(n1826), .Z(n823) );
  NR3SVTX6 U338 ( .A(n772), .B(n696), .C(n571), .Z(n845) );
  IVSVTX10 U339 ( .A(m1[13]), .Z(n920) );
  ND3SVTX4 U340 ( .A(n854), .B(n526), .C(n853), .Z(n44) );
  CTIVSVTX2 U341 ( .A(m1[0]), .Z(n843) );
  IVSVTX4 U342 ( .A(n1836), .Z(n970) );
  IVSVTX8 U343 ( .A(n702), .Z(n496) );
  ND2ASVTX6 U344 ( .A(n706), .B(n493), .Z(n743) );
  CTIVSVTX4 U345 ( .A(m1[1]), .Z(n853) );
  IVSVTX6 U346 ( .A(n677), .Z(n493) );
  IVSVTX10 U347 ( .A(m1[11]), .Z(n526) );
  IVSVTX10 U348 ( .A(n390), .Z(n391) );
  AO6SVTX2 U349 ( .A(n2009), .B(n703), .C(n1366), .Z(n1367) );
  AO7SVTX4 U350 ( .A(n1433), .B(n1432), .C(n981), .Z(n983) );
  F_ENSVTX2 U351 ( .A(n1816), .B(n1815), .Z(n1817) );
  F_ENSVTX2 U352 ( .A(n1389), .B(n1388), .Z(n1390) );
  AO6ABSVTX4 U353 ( .A(n128), .B(n1377), .C(n1376), .Z(n1385) );
  ENSVTX8 U354 ( .A(n1968), .B(n1967), .Z(m2[15]) );
  IVSVTX4 U355 ( .A(n1966), .Z(n1967) );
  AO7SVTX6 U356 ( .A(n1719), .B(n1722), .C(n1721), .Z(n1771) );
  F_EOSVTX2 U357 ( .A(n2039), .B(n2038), .Z(n2040) );
  AO6SVTX2 U358 ( .A(n102), .B(n2037), .C(n2036), .Z(n2038) );
  F_ENSVTX2 U359 ( .A(n1917), .B(n1916), .Z(n1926) );
  NR2SVTX2 U360 ( .A(n2013), .B(n2018), .Z(n2014) );
  F_ENSVTX2 U361 ( .A(n1357), .B(n1356), .Z(n1377) );
  F_ENSVTX2 U362 ( .A(n1702), .B(n1701), .Z(n1703) );
  F_ENSVTX2 U363 ( .A(n1666), .B(n1665), .Z(n1667) );
  AO6SVTX2 U364 ( .A(n1892), .B(n1890), .C(n1891), .Z(n1665) );
  AO3SVTX6 U365 ( .A(n128), .B(n1606), .C(n1605), .D(n1604), .Z(m2[7]) );
  AO6SVTX2 U366 ( .A(n1595), .B(n806), .C(n1594), .Z(n1596) );
  IVSVTX2 U367 ( .A(n1593), .Z(n1594) );
  AO6SVTX2 U368 ( .A(n1776), .B(n1775), .C(n1774), .Z(n1777) );
  AO2SVTX2 U369 ( .A(n673), .B(n1692), .C(n543), .D(n1691), .Z(n1698) );
  EOSVTX2 U370 ( .A(n1687), .B(n1686), .Z(n1692) );
  ND4SVTX6 U371 ( .A(n1736), .B(n1735), .C(n1734), .D(n1733), .Z(m2[4]) );
  ND2SVTX2 U372 ( .A(n1703), .B(n673), .Z(n1736) );
  AN3CSVTX4 U373 ( .A(n1994), .B(n1992), .C(n693), .Z(n2000) );
  F_ENSVTX2 U374 ( .A(n1423), .B(n1422), .Z(n1425) );
  AO7SVTX2 U375 ( .A(n1421), .B(n1813), .C(n1420), .Z(n1422) );
  ND4SVTX6 U376 ( .A(n1676), .B(n1675), .C(n1674), .D(n1673), .Z(m2[3]) );
  ND2SVTX2 U377 ( .A(n1667), .B(n673), .Z(n1675) );
  AO6SVTX2 U378 ( .A(n1951), .B(n806), .C(n1950), .Z(n1960) );
  ND2SVTX2 U379 ( .A(n1949), .B(n529), .Z(n1950) );
  F_EOSVTX2 U380 ( .A(n1368), .B(n1367), .Z(n1369) );
  ND3ABSVTX6 U381 ( .A(n640), .B(n639), .C(n638), .Z(m2[14]) );
  ND4SVTX6 U382 ( .A(n1430), .B(n1429), .C(n1428), .D(n1427), .Z(m2[10]) );
  EOSVTX2 U383 ( .A(n1764), .B(n1763), .Z(n1765) );
  AO7SVTX4 U384 ( .A(n1584), .B(n1701), .C(n1583), .Z(n1739) );
  ND2ASVTX8 U385 ( .A(n388), .B(n387), .Z(n1978) );
  NR3SVTX4 U386 ( .A(n2013), .B(n824), .C(n1325), .Z(n267) );
  F_EOSVTX2 U387 ( .A(n1956), .B(n1955), .Z(n1957) );
  ND3SVTX4 U388 ( .A(n777), .B(n970), .C(n393), .Z(n480) );
  ND2SVTX2 U389 ( .A(n777), .B(n504), .Z(n503) );
  AO7ASVTX6 U390 ( .A(n777), .B(n6), .C(m1[13]), .Z(n5) );
  ENSVTX2 U391 ( .A(n1445), .B(n1444), .Z(n1446) );
  ND4SVTX6 U392 ( .A(n1474), .B(n1473), .C(n1472), .D(n1471), .Z(m2[5]) );
  AO3SVTX6 U393 ( .A(n1424), .B(n747), .C(n1349), .D(n1348), .Z(m2[12]) );
  ENSVTX8 U394 ( .A(n155), .B(n1649), .Z(m2[18]) );
  AO7SVTX6 U395 ( .A(n1977), .B(n197), .C(n724), .Z(n1649) );
  AO2SVTX2 U396 ( .A(n1426), .B(n678), .C(n1425), .D(n1718), .Z(n1427) );
  NR2SVTX2 U397 ( .A(m1[6]), .B(n1628), .Z(n1773) );
  IVSVTX8 U398 ( .A(n412), .Z(n1531) );
  CTBUFSVTX4 U399 ( .A(n327), .Z(n189) );
  IVSVTX8 U400 ( .A(n1352), .Z(n339) );
  NR2SVTX4 U401 ( .A(n1264), .B(n1), .Z(n1165) );
  IVSVTX4 U402 ( .A(m1[16]), .Z(n919) );
  IVSVTX12 U403 ( .A(m1[19]), .Z(n869) );
  ND2SVTX4 U404 ( .A(n607), .B(n1453), .Z(n380) );
  NR2SVTX4 U405 ( .A(n381), .B(n682), .Z(n1453) );
  ND3ASVTX8 U406 ( .A(n1948), .B(n529), .C(n1958), .Z(n483) );
  AO7SVTX8 U407 ( .A(n1693), .B(n1895), .C(n1896), .Z(n35) );
  NR2SVTX4 U408 ( .A(n823), .B(n817), .Z(n17) );
  NR2SVTX4 U409 ( .A(n4), .B(n3), .Z(n1281) );
  ND2SVTX4 U410 ( .A(n1278), .B(n181), .Z(n3) );
  NR2SVTX4 U411 ( .A(n1280), .B(n1279), .Z(n4) );
  AO6SVTX6 U412 ( .A(n532), .B(n1226), .C(n738), .Z(n193) );
  ND2ASVTX8 U413 ( .A(n952), .B(n216), .Z(n1387) );
  ND2SVTX4 U414 ( .A(n5), .B(n1824), .Z(n952) );
  IVSVTX4 U415 ( .A(n493), .Z(n6) );
  AO7ABSVTX8 U416 ( .A(n728), .B(n133), .C(n1139), .Z(n450) );
  ND2SVTX8 U417 ( .A(n813), .B(n274), .Z(n814) );
  NR2SVTX4 U418 ( .A(n1230), .B(n1229), .Z(n1232) );
  ND2ASVTX8 U419 ( .A(n310), .B(n309), .Z(n311) );
  IVSVTX10 U420 ( .A(n390), .Z(n699) );
  ENSVTX8 U421 ( .A(n761), .B(n329), .Z(n214) );
  BFSVTX1 U422 ( .A(m1[23]), .Z(n11) );
  IVSVTX4 U423 ( .A(n81), .Z(n678) );
  IVSVTX6 U424 ( .A(n1083), .Z(n397) );
  AO6SVTX8 U425 ( .A(n922), .B(n1688), .C(n921), .Z(n1459) );
  IVSVTX8 U426 ( .A(n279), .Z(n282) );
  IVSVTX8 U427 ( .A(m1[9]), .Z(n828) );
  IVSVTX10 U428 ( .A(n705), .Z(n706) );
  AO7SVTX6 U429 ( .A(n528), .B(n625), .C(n658), .Z(n568) );
  AO7SVTX8 U430 ( .A(n81), .B(n252), .C(n251), .Z(n625) );
  IVSVTX8 U431 ( .A(n2031), .Z(n314) );
  NR2SVTX8 U432 ( .A(n628), .B(n561), .Z(n1992) );
  ND2ASVTX8 U433 ( .A(n171), .B(n709), .Z(n888) );
  BFSVTX4 U434 ( .A(m1[18]), .Z(n12) );
  ND2ASVTX8 U435 ( .A(n14), .B(n463), .Z(n462) );
  IVSVTX4 U436 ( .A(n845), .Z(n183) );
  AO6SVTX8 U437 ( .A(n1320), .B(n1157), .C(n1156), .Z(n29) );
  ND2ASVTX4 U438 ( .A(n1500), .B(n889), .Z(n774) );
  ND2ASVTX8 U439 ( .A(n15), .B(n407), .Z(n406) );
  ND2ASVTX8 U440 ( .A(n204), .B(n467), .Z(n1279) );
  IVSVTX4 U441 ( .A(n16), .Z(n269) );
  ND3SVTX6 U442 ( .A(n66), .B(n220), .C(n17), .Z(n16) );
  AO7ABSVTX4 U443 ( .A(n950), .B(n918), .C(n917), .Z(n587) );
  IVSVTX8 U444 ( .A(n391), .Z(n352) );
  BFSVTX1 U445 ( .A(n1353), .Z(n18) );
  NR3SVTX8 U446 ( .A(n427), .B(n224), .C(n223), .Z(n443) );
  AO7SVTX6 U447 ( .A(n887), .B(n443), .C(n488), .Z(n146) );
  ND3ASVTX8 U448 ( .A(n710), .B(n226), .C(n83), .Z(n560) );
  IVSVTX12 U449 ( .A(m1[11]), .Z(n813) );
  AO7SVTX6 U450 ( .A(n982), .B(n983), .C(n1431), .Z(n1582) );
  ND2SVTX4 U451 ( .A(n1433), .B(n1432), .Z(n1431) );
  ND2SVTX4 U452 ( .A(m1[2]), .B(n353), .Z(n1693) );
  AO7SVTX6 U453 ( .A(n497), .B(n501), .C(n500), .Z(n520) );
  AN2SVTX8 U454 ( .A(n80), .B(n630), .Z(n501) );
  ND2SVTX4 U455 ( .A(n355), .B(n19), .Z(n2004) );
  ENSVTX8 U456 ( .A(n243), .B(n20), .Z(n239) );
  AO6SVTX8 U457 ( .A(n1008), .B(n1486), .C(n1485), .Z(n20) );
  IVSVTX10 U458 ( .A(m1[6]), .Z(n527) );
  BFSVTX6 U459 ( .A(n1548), .Z(n22) );
  ND2SVTX4 U460 ( .A(n496), .B(n966), .Z(n1705) );
  NR2SVTX4 U461 ( .A(n25), .B(n1045), .Z(n84) );
  ND2SVTX4 U462 ( .A(n175), .B(n1304), .Z(n26) );
  AO2SVTX6 U463 ( .A(n1290), .B(n1109), .C(n730), .D(n1494), .Z(n1291) );
  ND2ASVTX8 U464 ( .A(n1108), .B(n1496), .Z(n1111) );
  IVSVTX2 U465 ( .A(n1111), .Z(n1110) );
  ND2ASVTX8 U466 ( .A(n28), .B(n27), .Z(n1981) );
  IVSVTX4 U467 ( .A(n838), .Z(n27) );
  IVSVTX4 U468 ( .A(n950), .Z(n28) );
  F_EOSVTX2 U469 ( .A(n1159), .B(n29), .Z(n1160) );
  IVSVTX2 U470 ( .A(n1258), .Z(n1154) );
  IVSVTX8 U471 ( .A(m1[16]), .Z(n277) );
  ND2SVTX6 U472 ( .A(n1190), .B(n1189), .Z(n141) );
  NR2SVTX4 U473 ( .A(n1878), .B(n1873), .Z(n922) );
  NR2SVTX4 U474 ( .A(n1836), .B(n966), .Z(n1878) );
  AO1ASVTX6 U475 ( .A(n1597), .B(n502), .C(n1178), .D(n1177), .Z(n1179) );
  AO7SVTX6 U476 ( .A(n1623), .B(n943), .C(n1622), .Z(n1825) );
  IVSVTX4 U477 ( .A(n493), .Z(n30) );
  IVSVTX4 U478 ( .A(n706), .Z(n31) );
  ND4SVTX6 U479 ( .A(n806), .B(n1499), .C(n595), .D(n597), .Z(n594) );
  AO6CSVTX8 U480 ( .A(n311), .B(n367), .C(n1495), .Z(n366) );
  IVSVTX12 U481 ( .A(n353), .Z(n696) );
  IVSVTX6 U482 ( .A(n1884), .Z(n855) );
  NR3SVTX8 U483 ( .A(n34), .B(n238), .C(n33), .Z(n248) );
  ND2SVTX4 U484 ( .A(n237), .B(n236), .Z(n33) );
  IVSVTX12 U485 ( .A(m1[5]), .Z(n353) );
  AO6ASVTX8 U486 ( .A(n382), .B(n1694), .C(n35), .Z(n1452) );
  AO6SVTX4 U487 ( .A(n74), .B(n1504), .C(n1503), .Z(n598) );
  ND2SVTX4 U488 ( .A(n1539), .B(n22), .Z(n1537) );
  IVSVTX10 U489 ( .A(n795), .Z(n695) );
  AO6SVTX4 U490 ( .A(n74), .B(n1504), .C(n1520), .Z(n1521) );
  IVSVTX4 U491 ( .A(n503), .Z(n754) );
  ND4SVTX8 U492 ( .A(n393), .B(n739), .C(n277), .D(n754), .Z(n785) );
  IVSVTX10 U493 ( .A(n705), .Z(n701) );
  AO7SVTX6 U494 ( .A(n768), .B(n141), .C(n38), .Z(n1192) );
  IVSVTX4 U495 ( .A(n708), .Z(n38) );
  ND2SVTX4 U496 ( .A(n766), .B(n94), .Z(n708) );
  ND4ABSVTX8 U497 ( .A(n293), .B(n294), .C(n39), .D(n659), .Z(n354) );
  ND2SVTX4 U498 ( .A(n1540), .B(n1539), .Z(n721) );
  ND2SVTX6 U499 ( .A(n1488), .B(n1044), .Z(n1065) );
  BFSVTX12 U500 ( .A(n828), .Z(n162) );
  ND2SVTX6 U501 ( .A(n186), .B(n185), .Z(n1576) );
  AO6CSVTX8 U502 ( .A(n1805), .B(n1803), .C(n1802), .Z(n1413) );
  IVSVTX8 U503 ( .A(n1413), .Z(n516) );
  BFSVTX1 U504 ( .A(n1878), .Z(n40) );
  AO7SVTX8 U505 ( .A(n901), .B(n900), .C(n1811), .Z(n378) );
  IVSVTX6 U506 ( .A(n997), .Z(n1510) );
  IVSVTX4 U507 ( .A(n71), .Z(n41) );
  ND2ASVTX8 U508 ( .A(n41), .B(n214), .Z(n251) );
  ENSVTX8 U509 ( .A(n11), .B(n307), .Z(n303) );
  ND3SVTX8 U510 ( .A(n614), .B(n615), .C(n613), .Z(n1645) );
  AO6SVTX8 U511 ( .A(n1825), .B(n43), .C(n815), .Z(n2021) );
  IVSVTX4 U512 ( .A(n822), .Z(n43) );
  ND2SVTX4 U513 ( .A(n1404), .B(n814), .Z(n822) );
  IVSVTX8 U514 ( .A(n80), .Z(n77) );
  IVSVTX8 U515 ( .A(n2029), .Z(n181) );
  IVSVTX6 U516 ( .A(n326), .Z(n322) );
  NR2SVTX4 U517 ( .A(n44), .B(n91), .Z(n318) );
  AO7SVTX8 U518 ( .A(n1767), .B(n414), .C(n1768), .Z(n923) );
  BFSVTX1 U519 ( .A(n1738), .Z(n45) );
  BFSVTX1 U520 ( .A(n743), .Z(n46) );
  AO17SVTX6 U521 ( .A(n51), .B(n50), .C(n49), .D(n48), .Z(n834) );
  IVSVTX4 U522 ( .A(n935), .Z(n49) );
  IVSVTX4 U523 ( .A(n936), .Z(n50) );
  IVSVTX4 U524 ( .A(n1527), .Z(n51) );
  NR2SVTX4 U525 ( .A(m1[3]), .B(n966), .Z(n1865) );
  NR3SVTX8 U526 ( .A(n822), .B(n1327), .C(n1463), .Z(n220) );
  BFSVTX1 U527 ( .A(n1437), .Z(n52) );
  NR2SVTX2 U528 ( .A(n1185), .B(n1301), .Z(n1276) );
  IVSVTX4 U529 ( .A(n1287), .Z(n1289) );
  BFSVTX2 U530 ( .A(n2021), .Z(n188) );
  ND2SVTX4 U531 ( .A(n769), .B(n54), .Z(n1178) );
  NR2ASVTX6 U532 ( .A(n1516), .B(n714), .Z(n1164) );
  AN2SVTX4 U533 ( .A(n813), .B(n828), .Z(n943) );
  AO6SVTX8 U534 ( .A(n1995), .B(n562), .C(n55), .Z(n524) );
  AO7SVTX8 U535 ( .A(n1990), .B(n1217), .C(n1215), .Z(n55) );
  AO7SVTX4 U536 ( .A(n1353), .B(n628), .C(n1350), .Z(n56) );
  AO6CSVTX8 U537 ( .A(n74), .B(n1028), .C(n206), .Z(n1029) );
  IVSVTX4 U538 ( .A(n1115), .Z(n1026) );
  ND2SVTX4 U539 ( .A(m1[13]), .B(m1[16]), .Z(n1336) );
  ND2SVTX4 U540 ( .A(n493), .B(n58), .Z(n1811) );
  AO7SVTX8 U541 ( .A(n719), .B(n1272), .C(n440), .Z(n439) );
  BFSVTX1 U542 ( .A(n1771), .Z(n59) );
  BFSVTX1 U543 ( .A(n1434), .Z(n60) );
  ND3SVTX8 U544 ( .A(n348), .B(n346), .C(n347), .Z(n997) );
  ND3ABSVTX4 U545 ( .A(n1060), .B(n593), .C(n424), .Z(n427) );
  ND2SVTX2 U546 ( .A(n106), .B(n632), .Z(n1277) );
  AO7SVTX2 U547 ( .A(n1557), .B(n790), .C(n1519), .Z(n1520) );
  AN2SVTX0H U548 ( .A(n104), .B(n1256), .Z(n751) );
  IVSVTX2 U549 ( .A(n1096), .Z(n591) );
  IVSVTX0H U550 ( .A(n129), .Z(n163) );
  F_ND2SVTX0H U551 ( .A(n1359), .B(n21), .Z(n1363) );
  NR2SVTX0H U552 ( .A(n2035), .B(n1378), .Z(n2037) );
  IVSVTX0H U553 ( .A(n1706), .Z(n1707) );
  AO7SVTX6 U554 ( .A(n1797), .B(n1795), .C(n1796), .Z(n1912) );
  IVSVTX0H U555 ( .A(n1378), .Z(n1380) );
  F_ND2SVTX0H U556 ( .A(n2003), .B(n2002), .Z(n2011) );
  IVSVTX2 U557 ( .A(n848), .Z(n86) );
  B_ND2SVTX0H U558 ( .A(n1896), .B(n894), .Z(n1900) );
  F_ND2SVTX0H U559 ( .A(n1755), .B(n734), .Z(n1764) );
  IVSVTX0H U560 ( .A(n1929), .Z(n1316) );
  EOSVTX0H U561 ( .A(n1753), .B(n1752), .Z(n1766) );
  AO6SVTX1 U562 ( .A(n1924), .B(n806), .C(n745), .Z(n1925) );
  F_ND2SVTX0H U563 ( .A(n1488), .B(n1670), .Z(n1674) );
  F_ND2SVTX0H U564 ( .A(n678), .B(n1603), .Z(n1604) );
  OR2SVTX1 U565 ( .A(n757), .B(n1523), .Z(n61) );
  IVSVTX2 U566 ( .A(n599), .Z(n1078) );
  F_AN2SVTX2 U567 ( .A(n119), .B(n728), .Z(n62) );
  IVSVTX10 U568 ( .A(m1[13]), .Z(n274) );
  IVSVTX6 U569 ( .A(m1[13]), .Z(n507) );
  ND2SVTX2 U570 ( .A(m1[3]), .B(m1[1]), .Z(n819) );
  IVSVTX12 U571 ( .A(m1[3]), .Z(n854) );
  IVSVTX6 U572 ( .A(m1[3]), .Z(n657) );
  F_IVSVTX0H U573 ( .A(n23), .Z(n1757) );
  IVSVTX10 U574 ( .A(m1[23]), .Z(n791) );
  IVSVTX12 U575 ( .A(n950), .Z(n588) );
  BFSVTX12 U576 ( .A(n80), .Z(n143) );
  AO7NSVTX8 U577 ( .A(n1741), .B(n1747), .C(n1743), .Z(n63) );
  AO5SVTX4 U578 ( .A(n133), .B(n168), .C(n916), .Z(n177) );
  AO7SVTX4 U579 ( .A(n133), .B(n917), .C(n600), .Z(n64) );
  F_ND2SVTX0H U580 ( .A(n1114), .B(n1113), .Z(n65) );
  F_ND2ASVTX2 U581 ( .A(n813), .B(n355), .Z(n1417) );
  AN3SVTX6 U582 ( .A(n1326), .B(n1323), .C(n333), .Z(n66) );
  AO6ASVTX8 U583 ( .A(n1929), .B(n1314), .C(n392), .Z(n2034) );
  F_AN2SVTX2 U584 ( .A(n1525), .B(n1008), .Z(n67) );
  AO6NSVTX4 U585 ( .A(n102), .B(n1253), .C(n1254), .Z(n68) );
  ND2SVTX2 U586 ( .A(n76), .B(n728), .Z(n573) );
  AN3SVTX6 U587 ( .A(n1095), .B(n573), .C(n718), .Z(n69) );
  F_AN2SVTX2 U588 ( .A(n200), .B(n226), .Z(n70) );
  IVSVTX6 U589 ( .A(n366), .Z(n1526) );
  NR3ABSVTX2 U590 ( .A(n200), .B(n1119), .C(n1194), .Z(n1092) );
  ND2SVTX2 U591 ( .A(n113), .B(n1128), .Z(n1131) );
  ND2SVTX4 U592 ( .A(n933), .B(n136), .Z(n1128) );
  AO17SVTX6 U593 ( .A(n1810), .B(n378), .C(n605), .D(n1417), .Z(n377) );
  AO7SVTX6 U594 ( .A(n1738), .B(n1578), .C(n1579), .Z(n495) );
  IVSVTX8 U595 ( .A(m1[9]), .Z(n963) );
  ENSVTX8 U596 ( .A(n760), .B(n1043), .Z(n1044) );
  AO3SVTX8 U597 ( .A(n930), .B(n1365), .C(n406), .D(n2003), .Z(n1953) );
  ND2SVTX4 U598 ( .A(n246), .B(n107), .Z(n883) );
  IVSVTX4 U599 ( .A(n1342), .Z(n737) );
  IVSVTX12 U600 ( .A(m1[2]), .Z(n895) );
  AO6SVTX8 U601 ( .A(n1953), .B(n932), .C(n931), .Z(n409) );
  BFSVTX12 U602 ( .A(n706), .Z(n1592) );
  AO4SVTX4 U603 ( .A(n977), .B(n978), .C(n1664), .D(n1663), .Z(n975) );
  ND3ABSVTX6 U604 ( .A(m1[23]), .B(m1[20]), .C(n838), .Z(n891) );
  ND3SVTX4 U605 ( .A(n920), .B(n473), .C(n816), .Z(n786) );
  IVSVTX8 U606 ( .A(m1[4]), .Z(n390) );
  AO17CSVTX4 U607 ( .A(n1490), .B(n466), .C(n609), .D(n673), .Z(n1491) );
  IVSVTX8 U608 ( .A(n398), .Z(n608) );
  NR2ASVTX1 U609 ( .A(n1662), .B(n60), .Z(n1666) );
  BFSVTX4 U610 ( .A(n1653), .Z(n421) );
  AO6SVTX8 U611 ( .A(n452), .B(n232), .C(n450), .Z(n416) );
  AN2BSVTX8 U612 ( .A(n527), .B(m1[3]), .Z(n1873) );
  AO7SVTX8 U613 ( .A(n612), .B(n610), .C(n617), .Z(n616) );
  F_ND2SVTX1 U614 ( .A(n2004), .B(n2005), .Z(n1368) );
  AO7SVTX6 U615 ( .A(n1570), .B(n360), .C(n1574), .Z(n1577) );
  IVSVTX6 U616 ( .A(n1571), .Z(n1570) );
  IVSVTX8 U617 ( .A(n282), .Z(n1516) );
  AO6ASVTX8 U618 ( .A(n2033), .B(n2030), .C(n314), .Z(n343) );
  AO6SVTX8 U619 ( .A(n1758), .B(n862), .C(n861), .Z(n170) );
  AO7SVTX8 U620 ( .A(n1754), .B(n1759), .C(n1755), .Z(n861) );
  ND2SVTX2 U621 ( .A(n827), .B(n963), .Z(n826) );
  F_ND2ASVTX2 U622 ( .A(m1[10]), .B(n827), .Z(n727) );
  IVSVTX8 U623 ( .A(n827), .Z(n630) );
  IVSVTX8 U624 ( .A(n827), .Z(n1779) );
  IVSVTX8 U625 ( .A(n827), .Z(n702) );
  ND2SVTX4 U626 ( .A(n909), .B(n869), .Z(n559) );
  AO3CDSVTX1 U627 ( .A(n1557), .B(n990), .C(n1555), .D(n1556), .Z(n1558) );
  AO7SVTX4 U628 ( .A(n998), .B(n1557), .C(n1501), .Z(n912) );
  AO7SVTX8 U629 ( .A(n1266), .B(n666), .C(n1262), .Z(n1174) );
  IVSVTX6 U630 ( .A(n1263), .Z(n666) );
  IVSVTX12 U631 ( .A(n572), .Z(n593) );
  ND2ASVTX8 U632 ( .A(n403), .B(n550), .Z(n546) );
  ND4ABSVTX8 U633 ( .A(n242), .B(n240), .C(n244), .D(n234), .Z(n369) );
  AO7SVTX6 U634 ( .A(n127), .B(n126), .C(n1534), .Z(n294) );
  NR2SVTX2 U635 ( .A(n660), .B(n345), .Z(n556) );
  ND2SVTX4 U636 ( .A(n1209), .B(n71), .Z(n529) );
  AO6CSVTX8 U637 ( .A(n1654), .B(n421), .C(n420), .Z(n1655) );
  IVSVTX8 U638 ( .A(n526), .Z(n947) );
  NR2ASVTX6 U639 ( .A(n904), .B(n110), .Z(n672) );
  ND2SVTX4 U640 ( .A(n402), .B(n398), .Z(n423) );
  AO6SVTX8 U641 ( .A(n516), .B(n361), .C(n850), .Z(n1152) );
  NR2SVTX2 U642 ( .A(m1[12]), .B(m1[10]), .Z(n445) );
  ND3SVTX4 U643 ( .A(n462), .B(n530), .C(n1119), .Z(n71) );
  IVSVTX8 U644 ( .A(n299), .Z(n232) );
  BFSVTX12 U645 ( .A(n232), .Z(n1718) );
  IVSVTX2 U646 ( .A(n1573), .Z(n205) );
  AO7SVTX4 U647 ( .A(n603), .B(n550), .C(n256), .Z(n255) );
  AO6SVTX8 U648 ( .A(n1771), .B(n541), .C(n923), .Z(n924) );
  AO2SVTX6 U649 ( .A(n438), .B(n95), .C(n435), .D(n675), .Z(n615) );
  IVSVTX6 U650 ( .A(n626), .Z(n395) );
  IVSVTX10 U651 ( .A(n1505), .Z(n72) );
  IVSVTX8 U652 ( .A(n72), .Z(n73) );
  IVSVTX12 U653 ( .A(n72), .Z(n74) );
  ND2SVTX2 U654 ( .A(n678), .B(n1711), .Z(n1735) );
  NR2ASVTX2 U655 ( .A(n1295), .B(n1294), .Z(n1296) );
  ND2SVTX2 U656 ( .A(n1108), .B(n1109), .Z(n578) );
  CTIVSVTX2 U657 ( .A(n1010), .Z(n1532) );
  IVSVTX2 U658 ( .A(n1492), .Z(n78) );
  CTIVSVTX2 U659 ( .A(n986), .Z(n542) );
  IVSVTX2 U660 ( .A(n729), .Z(n714) );
  OR2SVTX2 U661 ( .A(n2013), .B(n188), .Z(n375) );
  NR2SVTX2 U662 ( .A(n1494), .B(n730), .Z(n808) );
  CTIVSVTX2 U663 ( .A(n988), .Z(n794) );
  NR2SVTX2 U664 ( .A(n2006), .B(n700), .Z(n2008) );
  AO6SVTX4 U665 ( .A(n871), .B(n1041), .C(n870), .Z(n1484) );
  B_ND2SVTX1 U666 ( .A(n1935), .B(n1937), .Z(n1415) );
  OR2SVTX2 U667 ( .A(n1033), .B(n1032), .Z(n1034) );
  ND2SVTX2 U668 ( .A(n940), .B(n801), .Z(n1073) );
  IVSVTX6 U669 ( .A(n1171), .Z(n117) );
  B_ND2SVTX1 U670 ( .A(n1612), .B(n1613), .Z(n1618) );
  B_ND2SVTX1 U671 ( .A(n1637), .B(n1601), .Z(n1602) );
  ND2SVTX2 U672 ( .A(n933), .B(m1[25]), .Z(n1477) );
  CTIVSVTX6 U673 ( .A(n801), .Z(n75) );
  B_ND2SVTX1 U674 ( .A(n138), .B(n896), .Z(n1695) );
  IVSVTX4 U675 ( .A(n938), .Z(n94) );
  CTIVSVTX2 U676 ( .A(n1739), .Z(n1585) );
  AO7SVTX4 U677 ( .A(n437), .B(n68), .C(n436), .Z(n435) );
  CTIVSVTX2 U678 ( .A(n1187), .Z(n1184) );
  CTIVSVTX2 U679 ( .A(n1293), .Z(n1294) );
  CTIVSVTX2 U680 ( .A(n1145), .Z(n291) );
  MUX21NSVTX2 U681 ( .A(n1073), .B(n1144), .S(n1145), .Z(n290) );
  ND2SVTX6 U682 ( .A(n1144), .B(n101), .Z(n1185) );
  NR2SVTX2 U683 ( .A(n1136), .B(n1137), .Z(n513) );
  CTIVSVTX2 U684 ( .A(n631), .Z(n986) );
  ND2SVTX4 U685 ( .A(n1072), .B(n1071), .Z(n324) );
  CTIVSVTX4 U686 ( .A(n1497), .Z(n367) );
  IVSVTX2 U687 ( .A(n1106), .Z(n1108) );
  B_ND2SVTX1 U688 ( .A(n2012), .B(n148), .Z(n2024) );
  F_AN2SVTX2 U689 ( .A(n1122), .B(n1121), .Z(n1126) );
  CTIVSVTX2 U690 ( .A(n1173), .Z(n1170) );
  ND2SVTX4 U691 ( .A(n87), .B(n75), .Z(n1144) );
  CTIVSVTX2 U692 ( .A(n971), .Z(n196) );
  NR2SVTX2 U693 ( .A(n901), .B(n900), .Z(n1812) );
  B_ND2SVTX1 U694 ( .A(n1819), .B(n506), .Z(n1823) );
  B_ND2SVTX1 U695 ( .A(n166), .B(n1810), .Z(n1816) );
  CTIVSVTX2 U696 ( .A(n1932), .Z(n1933) );
  IVSVTX6 U697 ( .A(n277), .Z(n88) );
  IVSVTX0H U698 ( .A(n1935), .Z(n1936) );
  ND2SVTX6 U699 ( .A(n807), .B(n990), .Z(n250) );
  ND2SVTX2 U700 ( .A(n1013), .B(n1016), .Z(n488) );
  IVSVTX4 U701 ( .A(n117), .Z(n914) );
  IVSVTX2 U702 ( .A(n887), .Z(n565) );
  B_ND2SVTX2 U703 ( .A(n1017), .B(n773), .Z(n1199) );
  CTBUFSVTX2 U704 ( .A(n1454), .Z(n1746) );
  CTIVSVTX2 U705 ( .A(n893), .Z(n349) );
  IVSVTX2 U706 ( .A(n1845), .Z(n115) );
  B_ND2SVTX1 U707 ( .A(n1713), .B(n1714), .Z(n1671) );
  ND2SVTX6 U708 ( .A(n249), .B(n248), .Z(n1540) );
  B_ND2SVTX2 U709 ( .A(n1683), .B(n1488), .Z(n1699) );
  ND2ASVTX6 U710 ( .A(n99), .B(n673), .Z(n1096) );
  ND2SVTX2 U711 ( .A(n673), .B(n1446), .Z(n1474) );
  AO4SVTX1 U712 ( .A(n1829), .B(n718), .C(n1322), .D(n505), .Z(n1831) );
  AO17SVTX2 U713 ( .A(n1185), .B(n1187), .C(n1186), .D(n665), .Z(n758) );
  ND2SVTX4 U714 ( .A(n83), .B(n341), .Z(n938) );
  CTIVSVTX2 U715 ( .A(n1948), .Z(n1949) );
  IVSVTX8 U716 ( .A(n434), .Z(n2029) );
  F_EOSVTX2 U717 ( .A(n1163), .B(n1531), .Z(n502) );
  ND2SVTX2 U718 ( .A(n1187), .B(n1186), .Z(n665) );
  NR2ASVTX4 U719 ( .A(n434), .B(n290), .Z(n289) );
  NR3SVTX2 U720 ( .A(n914), .B(n1170), .C(n670), .Z(n336) );
  NR2SVTX4 U721 ( .A(n1497), .B(n1492), .Z(n1528) );
  B_ND2SVTX2 U722 ( .A(n603), .B(n555), .Z(n404) );
  NR2SVTX2 U723 ( .A(n1052), .B(n1051), .Z(n1050) );
  IVSVTX4 U724 ( .A(n1186), .Z(n204) );
  CTIVSVTX2 U725 ( .A(n1165), .Z(n670) );
  NR3SVTX2 U726 ( .A(n1018), .B(n1017), .C(n1016), .Z(n1020) );
  ND2SVTX2 U727 ( .A(n846), .B(n85), .Z(n1018) );
  IVSVTX2 U728 ( .A(n1954), .Z(n1271) );
  AO7SVTX4 U729 ( .A(n551), .B(n672), .C(n1270), .Z(n931) );
  ND2SVTX4 U730 ( .A(n85), .B(n432), .Z(n223) );
  B_ND2SVTX2 U731 ( .A(n1937), .B(n1933), .Z(n1939) );
  CTIVSVTX2 U732 ( .A(n1812), .Z(n1419) );
  CTIVSVTX2 U733 ( .A(n112), .Z(n263) );
  B_ND2SVTX2 U734 ( .A(n1417), .B(n1416), .Z(n1423) );
  CTIVSVTX2 U735 ( .A(n1011), .Z(n603) );
  IVSVTX0H U736 ( .A(n1810), .Z(n902) );
  CTIVSVTX2 U737 ( .A(n1161), .Z(n112) );
  IVSVTX2 U738 ( .A(n1210), .Z(n865) );
  NR4SVTX6 U739 ( .A(n696), .B(n455), .C(n460), .D(n203), .Z(n454) );
  NR2SVTX6 U740 ( .A(n731), .B(n1580), .Z(n964) );
  B_ND2SVTX2 U741 ( .A(n499), .B(n498), .Z(n980) );
  B_ND2SVTX1 U742 ( .A(n1588), .B(n151), .Z(n1589) );
  B_ND2SVTX1 U743 ( .A(n1875), .B(n1874), .Z(n1880) );
  NR2SVTX6 U744 ( .A(n920), .B(n475), .Z(n1360) );
  IVSVTX12 U745 ( .A(n904), .Z(n76) );
  B_ND2SVTX1 U746 ( .A(n1623), .B(n46), .Z(n1591) );
  IVSVTX8 U747 ( .A(m1[22]), .Z(n795) );
  CTIVSVTX2 U748 ( .A(n1975), .Z(n724) );
  ND2SVTX2 U749 ( .A(n1390), .B(n673), .Z(n1430) );
  ND3ASVTX6 U750 ( .A(n836), .B(n835), .C(n834), .Z(n939) );
  AO6SVTX2 U751 ( .A(n1994), .B(n1915), .C(n1912), .Z(n1388) );
  B_ND2SVTX2 U752 ( .A(n678), .B(n1640), .Z(n1641) );
  AO8SVTX2 U753 ( .A(n676), .B(n1355), .C(n1994), .D(n1354), .Z(n1356) );
  ND2SVTX4 U754 ( .A(n232), .B(n245), .Z(n244) );
  IVSVTX4 U755 ( .A(n95), .Z(n681) );
  B_ND2SVTX2 U756 ( .A(n95), .B(n1400), .Z(n1429) );
  CTBUFSVTX4 U757 ( .A(n230), .Z(n226) );
  ND2ASVTX6 U758 ( .A(n227), .B(n230), .Z(n228) );
  ND2SVTX6 U759 ( .A(n809), .B(n1165), .Z(n1492) );
  CTIVSVTX2 U760 ( .A(n285), .Z(n284) );
  ND4ABSVTX6 U761 ( .A(n119), .B(n86), .C(n671), .D(n847), .Z(n1242) );
  ND2SVTX4 U762 ( .A(n545), .B(n311), .Z(n1286) );
  AO1CDSVTX2 U763 ( .A(n276), .B(n1466), .C(n629), .D(n1465), .Z(n1785) );
  F_ND2ASVTX2 U764 ( .A(n1052), .B(n1049), .Z(n1059) );
  NR2ASVTX2 U765 ( .A(n1952), .B(n1271), .Z(n558) );
  IVSVTX2 U766 ( .A(n1143), .Z(n332) );
  ND2SVTX4 U767 ( .A(n788), .B(n787), .Z(n261) );
  ND2ASVTX6 U768 ( .A(n1142), .B(n1244), .Z(n331) );
  ND3SVTX6 U769 ( .A(n778), .B(n780), .C(n779), .Z(n1201) );
  B_ND2SVTX2 U770 ( .A(n1144), .B(n1073), .Z(n581) );
  ND2SVTX4 U771 ( .A(n787), .B(n788), .Z(n671) );
  IVSVTX6 U772 ( .A(n1482), .Z(n1280) );
  NR2SVTX6 U773 ( .A(n1072), .B(n1071), .Z(n1142) );
  AO6CSVTX6 U774 ( .A(n540), .B(n933), .C(n669), .Z(n788) );
  B_ND2SVTX1 U775 ( .A(n1270), .B(n1269), .Z(n759) );
  NR2SVTX4 U776 ( .A(n1127), .B(n1129), .Z(n1100) );
  CTIVSVTX2 U777 ( .A(n1325), .Z(n2016) );
  ND3SVTX4 U778 ( .A(n647), .B(n645), .C(n646), .Z(n1229) );
  ND2SVTX6 U779 ( .A(n749), .B(n1981), .Z(n868) );
  IVSVTX4 U780 ( .A(n1073), .Z(n1244) );
  AO6SVTX6 U781 ( .A(n749), .B(n866), .C(n865), .Z(n867) );
  CTIVSVTX4 U782 ( .A(n570), .Z(n2012) );
  IVSVTX6 U783 ( .A(n1222), .Z(n1795) );
  CTIVSVTX2 U784 ( .A(n1166), .Z(n286) );
  B_ND2SVTX2 U785 ( .A(n118), .B(n1907), .Z(n1908) );
  AN2SVTX4 U786 ( .A(n338), .B(n587), .Z(n655) );
  B_ND2SVTX1 U787 ( .A(n1615), .B(n1614), .Z(n1590) );
  IVSVTX8 U788 ( .A(n903), .Z(n1314) );
  B_ND2SVTX1 U789 ( .A(n115), .B(n1846), .Z(n1847) );
  AO7SVTX4 U790 ( .A(n1464), .B(n1727), .C(n1726), .Z(n831) );
  CTAN2BSVTX4 U791 ( .A(n807), .B(n933), .Z(n1104) );
  CTBUFSVTX4 U792 ( .A(n716), .Z(n136) );
  IVSVTX8 U793 ( .A(n355), .Z(n89) );
  F_AN2SVTX2 U794 ( .A(n1664), .B(n1663), .Z(n1891) );
  IVSVTX4 U795 ( .A(n485), .Z(n487) );
  IVSVTX2 U796 ( .A(n795), .Z(n431) );
  IVSVTX0H U797 ( .A(n896), .Z(n1898) );
  ND2SVTX4 U798 ( .A(m1[1]), .B(n854), .Z(n1841) );
  IVSVTX4 U799 ( .A(m1[1]), .Z(n139) );
  NR2SVTX6 U800 ( .A(n1191), .B(n1192), .Z(n1644) );
  F_ENSVTX2 U801 ( .A(n1801), .B(n1800), .Z(n1835) );
  AO7SVTX2 U802 ( .A(n149), .B(n1798), .C(n1797), .Z(n1800) );
  NR2SVTX2 U803 ( .A(n1999), .B(n2000), .Z(n642) );
  AO4SVTX2 U804 ( .A(n1322), .B(n920), .C(n718), .D(n1333), .Z(n1334) );
  AO4SVTX2 U805 ( .A(n1322), .B(n496), .C(n1789), .D(n718), .Z(n1790) );
  B_ND2SVTX2 U806 ( .A(n1894), .B(n673), .Z(n1903) );
  IVSVTX4 U807 ( .A(n218), .Z(n993) );
  NR3SVTX4 U808 ( .A(n106), .B(n1280), .C(n82), .Z(n557) );
  AO7SVTX2 U809 ( .A(n98), .B(n1292), .C(n1291), .Z(n1299) );
  AO4SVTX4 U810 ( .A(n403), .B(n1056), .C(n602), .D(n404), .Z(n254) );
  IVSVTX10 U811 ( .A(n82), .Z(n673) );
  ND2ASVTX4 U812 ( .A(n215), .B(n228), .Z(n218) );
  NR2SVTX6 U813 ( .A(n811), .B(n98), .Z(n935) );
  CTIVSVTX2 U814 ( .A(n693), .Z(n676) );
  IVSVTX4 U815 ( .A(n97), .Z(n83) );
  F_ENSVTX2 U816 ( .A(n1126), .B(n1125), .Z(n452) );
  NR2SVTX2 U817 ( .A(n1054), .B(n1053), .Z(n1055) );
  IVSVTX4 U818 ( .A(n1286), .Z(n98) );
  ND2ASVTX4 U819 ( .A(n117), .B(n1201), .Z(n385) );
  ND2SVTX4 U820 ( .A(n1100), .B(n84), .Z(n555) );
  IVSVTX4 U821 ( .A(n1237), .Z(n100) );
  IVSVTX4 U822 ( .A(n311), .Z(n1496) );
  B_ND2SVTX1 U823 ( .A(n1355), .B(n18), .Z(n1345) );
  IVSVTX2 U824 ( .A(n1074), .Z(n518) );
  AO6SVTX4 U825 ( .A(n311), .B(n1035), .C(n1105), .Z(n539) );
  CTIVSVTX2 U826 ( .A(n1176), .Z(n715) );
  IVSVTX4 U827 ( .A(n1142), .Z(n101) );
  NR2SVTX6 U828 ( .A(n868), .B(n1983), .Z(n1258) );
  AO7SVTX4 U829 ( .A(n1097), .B(n1047), .C(n1098), .Z(n1048) );
  B_ND2SVTX2 U830 ( .A(n1098), .B(n250), .Z(n1101) );
  IVSVTX2 U831 ( .A(n1019), .Z(n549) );
  ND2SVTX4 U832 ( .A(n830), .B(n266), .Z(n1329) );
  IVSVTX2 U833 ( .A(n1203), .Z(n1204) );
  F_AN2SVTX2 U834 ( .A(n1079), .B(n599), .Z(n1082) );
  IVSVTX2 U835 ( .A(n1041), .Z(n1006) );
  B_ND2SVTX2 U836 ( .A(n551), .B(n1952), .Z(n1956) );
  ND2ASVTX6 U837 ( .A(n1502), .B(n1287), .Z(n1497) );
  NR2SVTX2 U838 ( .A(n1266), .B(n1267), .Z(n618) );
  CTIVSVTX2 U839 ( .A(n1116), .Z(n1025) );
  IVSVTX4 U840 ( .A(n531), .Z(n1796) );
  AO7ABSVTX4 U841 ( .A(n559), .B(n810), .C(n1133), .Z(n310) );
  B_ND2SVTX2 U842 ( .A(n1262), .B(n1263), .Z(n1267) );
  CTIVSVTX4 U843 ( .A(n159), .Z(n1502) );
  IVSVTX2 U844 ( .A(n802), .Z(n803) );
  B_ND2SVTX2 U845 ( .A(n744), .B(n57), .Z(n1132) );
  IVSVTX4 U846 ( .A(n880), .Z(n85) );
  ND2SVTX4 U847 ( .A(n116), .B(n88), .Z(n2017) );
  ND4ABSVTX6 U848 ( .A(n571), .B(n696), .C(n459), .D(n844), .Z(n880) );
  B_ND2SVTX1 U849 ( .A(n1867), .B(n1866), .Z(n1872) );
  IVSVTX4 U850 ( .A(n838), .Z(n110) );
  B_ND2SVTX2 U851 ( .A(n1436), .B(n1435), .Z(n1890) );
  CTIVSVTX2 U852 ( .A(n1148), .Z(n1124) );
  CTIVSVTX2 U853 ( .A(n1477), .Z(n1011) );
  NR2SVTX4 U854 ( .A(m1[27]), .B(n893), .Z(n848) );
  IVSVTX0H U855 ( .A(n1609), .Z(n1588) );
  AO7SVTX2 U856 ( .A(n1784), .B(n1782), .C(n1780), .Z(n829) );
  NR2ASVTX4 U857 ( .A(n352), .B(n1837), .Z(n1845) );
  CTIVSVTX2 U858 ( .A(n881), .Z(n773) );
  IVSVTX4 U859 ( .A(m1[25]), .Z(n1529) );
  IVSVTX2 U860 ( .A(n501), .Z(n498) );
  IVSVTX10 U861 ( .A(m1[24]), .Z(n910) );
  IVSVTX10 U862 ( .A(n1830), .Z(n80) );
  ND3SVTX4 U863 ( .A(n1574), .B(n1572), .C(n187), .Z(n1575) );
  IVSVTX4 U864 ( .A(n423), .Z(n422) );
  CTIVSVTX2 U865 ( .A(n389), .Z(n388) );
  NR2SVTX2 U866 ( .A(n128), .B(n641), .Z(n640) );
  IVSVTX2 U867 ( .A(n1561), .Z(n93) );
  AO6SVTX2 U868 ( .A(n95), .B(n1633), .C(n1632), .Z(n1642) );
  AO6SVTX2 U869 ( .A(n1335), .B(n678), .C(n1334), .Z(n1349) );
  NR2SVTX6 U870 ( .A(n1193), .B(n1181), .Z(n1974) );
  IVSVTX4 U871 ( .A(n358), .Z(n347) );
  IVSVTX2 U872 ( .A(n1273), .Z(n564) );
  ND3SVTX4 U873 ( .A(n789), .B(n1528), .C(n368), .Z(n597) );
  AO7SVTX6 U874 ( .A(n8), .B(n368), .C(n578), .Z(n577) );
  IVSVTX6 U875 ( .A(n680), .Z(n1284) );
  F_ENSVTX2 U876 ( .A(n1587), .B(n1586), .Z(n1606) );
  F_ND2SVTX1 U877 ( .A(n1488), .B(n1450), .Z(n1473) );
  CTIVSVTX4 U878 ( .A(n1491), .Z(n242) );
  ND2ASVTX4 U879 ( .A(n1285), .B(n365), .Z(n1300) );
  ND3SVTX6 U880 ( .A(n137), .B(n1490), .C(n673), .Z(n241) );
  B_ND2SVTX2 U881 ( .A(n673), .B(n758), .Z(n768) );
  IVSVTX6 U882 ( .A(n365), .Z(n368) );
  AO6SVTX2 U883 ( .A(n1056), .B(n1479), .C(n1478), .Z(n1480) );
  IVSVTX2 U884 ( .A(n1103), .Z(n465) );
  IVSVTX2 U885 ( .A(n1276), .Z(n1283) );
  IVSVTX8 U886 ( .A(n634), .Z(n635) );
  NR3SVTX4 U887 ( .A(n2029), .B(n99), .C(n1102), .Z(n1103) );
  NR4ABSVTX4 U888 ( .A(n1302), .B(n804), .C(n2029), .D(n1301), .Z(n1303) );
  ND2ASVTX4 U889 ( .A(n78), .B(n1110), .Z(n576) );
  F_ND2ASVTX2 U890 ( .A(n393), .B(n225), .Z(n589) );
  B_ND2SVTX2 U891 ( .A(n543), .B(n1928), .Z(n161) );
  IVSVTX8 U892 ( .A(n210), .Z(n321) );
  IVSVTX4 U893 ( .A(n1528), .Z(n297) );
  CTBUFSVTX4 U894 ( .A(n728), .Z(n225) );
  ND2SVTX4 U895 ( .A(n539), .B(n538), .Z(n1037) );
  CTIVSVTX2 U896 ( .A(n1107), .Z(n124) );
  B_ND2SVTX2 U897 ( .A(n375), .B(n1370), .Z(n374) );
  F_ENSVTX2 U898 ( .A(n65), .B(n1117), .Z(n579) );
  CTBUFSVTX4 U899 ( .A(n1627), .Z(n165) );
  F_EOSVTX2 U900 ( .A(n1382), .B(n1381), .Z(n1383) );
  CTBUFSVTX4 U901 ( .A(n1167), .Z(n200) );
  AO4SVTX4 U902 ( .A(n1208), .B(n102), .C(n344), .D(n1203), .Z(n1205) );
  ND2SVTX2 U903 ( .A(n765), .B(n1202), .Z(n1948) );
  IVSVTX8 U904 ( .A(n228), .Z(n82) );
  CTBUFSVTX12 U905 ( .A(n698), .Z(n281) );
  IVSVTX4 U906 ( .A(n1076), .Z(n99) );
  IVSVTX0H U907 ( .A(n532), .Z(n142) );
  AO6SVTX2 U908 ( .A(n102), .B(n1380), .C(n1379), .Z(n1381) );
  B_ND2SVTX2 U909 ( .A(n1991), .B(n1990), .Z(n2001) );
  IVSVTX2 U910 ( .A(n558), .Z(n719) );
  ND2ASVTX4 U911 ( .A(n286), .B(n512), .Z(n285) );
  ND2ASVTX6 U912 ( .A(n1329), .B(n1328), .Z(n2015) );
  AO7NSVTX1 U913 ( .A(n2018), .B(n1370), .C(n2017), .Z(n2019) );
  ND2SVTX4 U914 ( .A(n976), .B(n984), .Z(n654) );
  NR3ABSVTX4 U915 ( .A(n911), .B(n447), .C(n884), .Z(n1515) );
  NR2SVTX6 U916 ( .A(n172), .B(n914), .Z(n227) );
  IVSVTX4 U917 ( .A(n864), .Z(n515) );
  AO7SVTX2 U918 ( .A(n1039), .B(n1006), .C(n1005), .Z(n1007) );
  ND2ASVTX4 U919 ( .A(n108), .B(n1174), .Z(n512) );
  AO6SVTX4 U920 ( .A(n736), .B(n775), .C(n774), .Z(n779) );
  F_ND2SVTX1 U921 ( .A(n1174), .B(n1173), .Z(n1175) );
  IVSVTX4 U922 ( .A(n1289), .Z(n545) );
  F_AN2SVTX2 U923 ( .A(n1501), .B(n999), .Z(n761) );
  AO7SVTX1 U924 ( .A(n1870), .B(n1869), .C(n1868), .Z(n1871) );
  AO7SVTX4 U925 ( .A(n1935), .B(n664), .C(n1931), .Z(n850) );
  B_ND2SVTX1 U926 ( .A(n1393), .B(n1819), .Z(n1397) );
  CTIVSVTX2 U927 ( .A(n1459), .Z(n1775) );
  F_AN2SVTX2 U928 ( .A(n1005), .B(n1040), .Z(n760) );
  IVSVTX4 U929 ( .A(n492), .Z(n1482) );
  ND3SVTX4 U930 ( .A(n105), .B(n511), .C(n892), .Z(n446) );
  IVSVTX2 U931 ( .A(n425), .Z(n846) );
  ND3SVTX4 U932 ( .A(n723), .B(n1811), .C(n1416), .Z(n383) );
  NR2SVTX6 U933 ( .A(n802), .B(n793), .Z(n492) );
  NR3SVTX4 U934 ( .A(n28), .B(n116), .C(n183), .Z(n468) );
  B_ND2SVTX1 U935 ( .A(n1931), .B(n849), .Z(n1941) );
  B_ND2SVTX1 U936 ( .A(n1324), .B(n1323), .Z(n1332) );
  B_ND2SVTX2 U937 ( .A(n1003), .B(n1002), .Z(n763) );
  B_ND2SVTX2 U938 ( .A(n1166), .B(n152), .Z(n1173) );
  IVSVTX0H U939 ( .A(n2013), .Z(n1371) );
  F_AN2SVTX2 U940 ( .A(n1907), .B(n1337), .Z(n703) );
  AO7SVTX1 U941 ( .A(n1898), .B(n1897), .C(n138), .Z(n1899) );
  B_ND2SVTX2 U942 ( .A(n1151), .B(n109), .Z(n1159) );
  IVSVTX4 U943 ( .A(n1249), .Z(n1252) );
  IVSVTX4 U944 ( .A(n898), .Z(n1416) );
  ND3SVTX4 U945 ( .A(n448), .B(n881), .C(n910), .Z(n470) );
  NR2SVTX1 U946 ( .A(n1770), .B(n164), .Z(n1776) );
  CTIVSVTX2 U947 ( .A(n1581), .Z(n1584) );
  IVSVTX4 U948 ( .A(n831), .Z(n150) );
  CTAN2BSVTX4 U949 ( .A(n669), .B(n1529), .Z(n1523) );
  CTIVSVTX2 U950 ( .A(n132), .Z(n1681) );
  IVSVTX2 U951 ( .A(n829), .Z(n830) );
  CTBUFSVTX12 U952 ( .A(n695), .Z(n168) );
  B_ND2SVTX1 U953 ( .A(n1852), .B(n1851), .Z(n1853) );
  IVSVTX4 U954 ( .A(n520), .Z(n519) );
  IVSVTX4 U955 ( .A(n940), .Z(n87) );
  B_ND2SVTX1 U956 ( .A(n1803), .B(n1802), .Z(n1809) );
  B_ND2SVTX2 U957 ( .A(n1712), .B(n376), .Z(n1716) );
  B_ND2SVTX1 U958 ( .A(n1784), .B(n1783), .Z(n1467) );
  F_ND2ASVTX2 U959 ( .A(n965), .B(n1442), .Z(n1443) );
  ND2ASVTX6 U960 ( .A(n657), .B(n153), .Z(n1884) );
  IVSVTX0H U961 ( .A(n1620), .Z(n1621) );
  IVSVTX4 U962 ( .A(n825), .Z(n1727) );
  CTIVSVTX6 U963 ( .A(n1607), .Z(n90) );
  IVSVTX8 U964 ( .A(n918), .Z(n91) );
  F_ND2SVTX0H U965 ( .A(m1[25]), .B(m1[24]), .Z(n1014) );
  IVSVTX6 U966 ( .A(n734), .Z(n1754) );
  CTBUFSVTX4 U967 ( .A(m1[24]), .Z(n1500) );
  IVSVTX2 U968 ( .A(n826), .Z(n1782) );
  IVSVTX4 U969 ( .A(n212), .Z(n160) );
  ND2SVTX2 U970 ( .A(n191), .B(n1307), .Z(n190) );
  IVSVTX2 U971 ( .A(n1308), .Z(n191) );
  ND3SVTX4 U972 ( .A(n161), .B(n1944), .C(n1927), .Z(m2[11]) );
  IVSVTX2 U973 ( .A(n169), .Z(n1650) );
  ND4SVTX4 U974 ( .A(n1864), .B(n1863), .C(n1862), .D(n1861), .Z(m2[0]) );
  ND4SVTX4 U975 ( .A(n1905), .B(n1904), .C(n1903), .D(n1902), .Z(m2[2]) );
  AO3ABSVTX4 U976 ( .A(n1718), .B(n1643), .C(n1642), .D(n1641), .Z(m2[8]) );
  ND4SVTX4 U977 ( .A(n1700), .B(n1699), .C(n1698), .D(n1697), .Z(m2[1]) );
  AO7NSVTX4 U978 ( .A(n128), .B(n1926), .C(n1925), .Z(n1927) );
  AO3SVTX4 U979 ( .A(n128), .B(n1794), .C(n1793), .D(n1792), .Z(m2[6]) );
  AO2SVTX2 U980 ( .A(n1364), .B(n678), .C(n165), .D(n89), .Z(n1375) );
  B_ND2SVTX2 U981 ( .A(n1889), .B(n678), .Z(n1904) );
  AO7ABSVTX2 U982 ( .A(n2042), .B(n678), .C(n2041), .Z(n639) );
  B_ND2SVTX2 U983 ( .A(n1844), .B(n678), .Z(n1863) );
  IVSVTX2 U984 ( .A(n2028), .Z(n638) );
  B_ND2SVTX2 U985 ( .A(n1718), .B(n1383), .Z(n1384) );
  B_ND2SVTX2 U986 ( .A(n1860), .B(n1718), .Z(n1861) );
  AO6SVTX2 U987 ( .A(n1832), .B(n543), .C(n1831), .Z(n1833) );
  ND3SVTX4 U988 ( .A(n1300), .B(n1299), .C(n1298), .Z(n175) );
  ND2ASVTX4 U989 ( .A(n996), .B(n995), .Z(n348) );
  B_ND2SVTX2 U990 ( .A(n1696), .B(n1718), .Z(n1697) );
  AO6SVTX2 U991 ( .A(n543), .B(n1732), .C(n1731), .Z(n1733) );
  B_ND2SVTX2 U992 ( .A(n1718), .B(n1457), .Z(n1472) );
  B_ND2SVTX2 U993 ( .A(n1718), .B(n1717), .Z(n1734) );
  IVSVTX2 U994 ( .A(n1506), .Z(n233) );
  ND2SVTX6 U995 ( .A(n1488), .B(n239), .Z(n231) );
  F_ENSVTX2 U996 ( .A(n1518), .B(n1480), .Z(n1481) );
  ND4SVTX6 U997 ( .A(n878), .B(n879), .C(n877), .D(n306), .Z(n305) );
  ND2SVTX4 U998 ( .A(n465), .B(n464), .Z(n400) );
  ND3SVTX4 U999 ( .A(n988), .B(n359), .C(n993), .Z(n835) );
  ND3ABSVTX6 U1000 ( .A(n1559), .B(n1021), .C(n342), .Z(n1194) );
  IVSVTX2 U1001 ( .A(n83), .Z(n679) );
  AO17SVTX6 U1002 ( .A(n297), .B(n910), .C(n1526), .D(n596), .Z(n595) );
  F_ENSVTX2 U1003 ( .A(n1034), .B(n1037), .Z(n1038) );
  AO8SVTX2 U1004 ( .A(n2015), .B(n2016), .C(n1371), .D(n374), .Z(n373) );
  NR2SVTX4 U1005 ( .A(n297), .B(n1527), .Z(n296) );
  F_AN2SVTX2 U1006 ( .A(n704), .B(n225), .Z(n745) );
  IVSVTX2 U1007 ( .A(n1195), .Z(n732) );
  AO7SVTX4 U1008 ( .A(n1559), .B(n1168), .C(n91), .Z(n769) );
  NR3ABSVTX6 U1009 ( .A(n1242), .B(n1241), .C(n1195), .Z(n342) );
  ND2ASVTX4 U1010 ( .A(n603), .B(n602), .Z(n256) );
  F_ENSVTX2 U1011 ( .A(n211), .B(n598), .Z(n245) );
  IVSVTX4 U1012 ( .A(n1627), .Z(n341) );
  IVSVTX4 U1013 ( .A(n262), .Z(n264) );
  IVSVTX8 U1014 ( .A(n1597), .Z(n95) );
  AO3SVTX1 U1015 ( .A(n188), .B(n2022), .C(n2020), .D(n2019), .Z(n2023) );
  AO7SVTX2 U1016 ( .A(n1786), .B(n1785), .C(n1784), .Z(n1787) );
  IVSVTX4 U1017 ( .A(n1242), .Z(n97) );
  ND2SVTX2 U1018 ( .A(n549), .B(n1020), .Z(n548) );
  IVSVTX2 U1019 ( .A(n530), .Z(n1021) );
  F_EOSVTX2 U1020 ( .A(n1716), .B(n1715), .Z(n1717) );
  ND4ABSVTX6 U1021 ( .A(n886), .B(n172), .C(n885), .D(n884), .Z(n530) );
  CTIVSVTX6 U1022 ( .A(n1231), .Z(n755) );
  NR2SVTX6 U1023 ( .A(n1219), .B(n1218), .Z(n656) );
  AO7SVTX4 U1024 ( .A(n694), .B(n489), .C(n349), .Z(n179) );
  ND3ABSVTX4 U1025 ( .A(n891), .B(n510), .C(n892), .Z(n1019) );
  ND2SVTX6 U1026 ( .A(n750), .B(n661), .Z(n1231) );
  IVSVTX6 U1027 ( .A(n604), .Z(n102) );
  ND2SVTX4 U1028 ( .A(n510), .B(n1133), .Z(n509) );
  ND2SVTX6 U1029 ( .A(n648), .B(n1662), .Z(n644) );
  NR2SVTX1 U1030 ( .A(n1920), .B(n1919), .Z(n1923) );
  B_ND2SVTX2 U1031 ( .A(n1361), .B(n1319), .Z(n1321) );
  AO7SVTX4 U1032 ( .A(n1251), .B(n1246), .C(n1248), .Z(n905) );
  B_ND2SVTX2 U1033 ( .A(n1266), .B(n1267), .Z(n1268) );
  IVSVTX4 U1034 ( .A(n247), .Z(n246) );
  ND2ASVTX6 U1035 ( .A(n1327), .B(n150), .Z(n266) );
  CTIVSVTX4 U1036 ( .A(n694), .Z(n103) );
  AO7SVTX4 U1037 ( .A(n1033), .B(n1036), .C(n1031), .Z(n1493) );
  AO7SVTX4 U1038 ( .A(n371), .B(n1918), .C(n1324), .Z(n812) );
  AO7SVTX4 U1039 ( .A(n1005), .B(n1001), .C(n1003), .Z(n870) );
  IVSVTX4 U1040 ( .A(n1387), .Z(n533) );
  IVSVTX2 U1041 ( .A(n486), .Z(n171) );
  AO3SVTX6 U1042 ( .A(n711), .B(n927), .C(n259), .D(n1392), .Z(n928) );
  AO7SVTX1 U1043 ( .A(n1748), .B(n156), .C(n1747), .Z(n1749) );
  B_ND2SVTX2 U1044 ( .A(n1885), .B(n1681), .Z(n1682) );
  B_ND2SVTX1 U1045 ( .A(n166), .B(n154), .Z(n1421) );
  B_ND2SVTX2 U1046 ( .A(n1148), .B(n1147), .Z(n1149) );
  B_ND2SVTX2 U1047 ( .A(n2033), .B(n2032), .Z(n1382) );
  OR2SVTX4 U1048 ( .A(n790), .B(n1477), .Z(n741) );
  B_ND2SVTX1 U1049 ( .A(n134), .B(n1458), .Z(n1461) );
  B_ND2SVTX2 U1050 ( .A(n1451), .B(n1747), .Z(n1456) );
  IVSVTX4 U1051 ( .A(n1255), .Z(n104) );
  AO7SVTX2 U1052 ( .A(n1772), .B(n164), .C(n134), .Z(n1774) );
  CTIVSVTX2 U1053 ( .A(n1123), .Z(n1147) );
  IVSVTX4 U1054 ( .A(n891), .Z(n105) );
  NR2SVTX1 U1055 ( .A(n1870), .B(n1677), .Z(n1679) );
  IVSVTX2 U1056 ( .A(n1489), .Z(n633) );
  IVSVTX4 U1057 ( .A(n804), .Z(n106) );
  B_ND2SVTX2 U1058 ( .A(n1841), .B(n1840), .Z(n1842) );
  NR2SVTX1 U1059 ( .A(n1745), .B(n156), .Z(n1750) );
  NR2SVTX6 U1060 ( .A(n1608), .B(n90), .Z(n900) );
  AO7NSVTX2 U1061 ( .A(n1843), .B(n753), .C(n1841), .Z(n771) );
  B_ND2SVTX2 U1062 ( .A(n1706), .B(n1708), .Z(n1669) );
  IVSVTX4 U1063 ( .A(n152), .Z(n108) );
  NR2SVTX1 U1064 ( .A(n1782), .B(n1781), .Z(n1788) );
  IVSVTX0H U1065 ( .A(n1405), .Z(n689) );
  AO7SVTX4 U1066 ( .A(n970), .B(n969), .C(n968), .Z(n1848) );
  IVSVTX2 U1067 ( .A(n1870), .Z(n157) );
  NR2SVTX4 U1068 ( .A(n1719), .B(n1658), .Z(n1769) );
  B_ND2SVTX2 U1069 ( .A(n1721), .B(n1720), .Z(n1725) );
  IVSVTX8 U1070 ( .A(n854), .Z(n772) );
  AO7SVTX6 U1071 ( .A(n1706), .B(n1704), .C(n1705), .Z(n1758) );
  CTIVSVTX4 U1072 ( .A(n1906), .Z(n118) );
  IVSVTX10 U1073 ( .A(m1[18]), .Z(n918) );
  IVSVTX2 U1074 ( .A(n1615), .Z(n712) );
  IVSVTX2 U1075 ( .A(n504), .Z(n477) );
  IVSVTX4 U1076 ( .A(n684), .Z(n1722) );
  IVSVTX4 U1077 ( .A(n720), .Z(n1704) );
  IVSVTX4 U1078 ( .A(n692), .Z(n1767) );
  IVSVTX10 U1079 ( .A(m1[10]), .Z(n1830) );
  AO3SVTX8 U1080 ( .A(n626), .B(n1553), .C(n1540), .D(n184), .Z(n360) );
  ND3ABSVTX6 U1081 ( .A(n680), .B(n528), .C(n623), .Z(n357) );
  ND3SVTX8 U1082 ( .A(n472), .B(n257), .C(n253), .Z(n528) );
  IVSVTX10 U1083 ( .A(n1498), .Z(n365) );
  ND2SVTX4 U1084 ( .A(n960), .B(n961), .Z(n1353) );
  EO3SVTX8 U1085 ( .A(m1[16]), .B(n475), .C(n683), .Z(n961) );
  ENSVTX8 U1086 ( .A(n1980), .B(n1979), .Z(m2[19]) );
  BFSVTX2 U1087 ( .A(n755), .Z(n122) );
  ND2SVTX4 U1088 ( .A(m1[6]), .B(n854), .Z(n894) );
  ND2ASVTX8 U1089 ( .A(n446), .B(n103), .Z(n884) );
  ND2SVTX4 U1090 ( .A(n916), .B(n915), .Z(n1031) );
  ND2SVTX4 U1091 ( .A(n115), .B(n196), .Z(n972) );
  IVSVTX8 U1092 ( .A(n91), .Z(n429) );
  IVSVTX8 U1093 ( .A(m1[12]), .Z(n777) );
  AO6SVTX8 U1094 ( .A(n1394), .B(n929), .C(n928), .Z(n411) );
  AO7SVTX4 U1095 ( .A(n1150), .B(n1256), .C(n1151), .Z(n514) );
  ND2SVTX4 U1096 ( .A(n260), .B(n1613), .Z(n713) );
  ND2SVTX4 U1097 ( .A(n123), .B(n704), .Z(n1613) );
  IVSVTX4 U1098 ( .A(n162), .Z(n123) );
  IVSVTX8 U1099 ( .A(n828), .Z(n1628) );
  IVSVTX12 U1100 ( .A(n1830), .Z(n677) );
  NR2SVTX4 U1101 ( .A(m1[9]), .B(n706), .Z(n504) );
  ND2ASVTX8 U1102 ( .A(n124), .B(n265), .Z(n575) );
  NR2SVTX4 U1103 ( .A(n296), .B(n1526), .Z(n127) );
  AO7CSVTX6 U1104 ( .A(n255), .B(n254), .C(n1597), .Z(n253) );
  AO7SVTX8 U1105 ( .A(n1876), .B(n1873), .C(n1875), .Z(n921) );
  F_AN2SVTX2 U1106 ( .A(n1024), .B(n1023), .Z(n752) );
  CTBUFSVTX8 U1107 ( .A(n411), .Z(n130) );
  NR2SVTX4 U1108 ( .A(n701), .B(n32), .Z(n1719) );
  ND3ASVTX8 U1109 ( .A(n442), .B(n179), .C(n146), .Z(n1119) );
  ND2SVTX4 U1110 ( .A(n2030), .B(n2032), .Z(n394) );
  ND2ASVTX8 U1111 ( .A(n131), .B(n957), .Z(n2030) );
  ND2SVTX4 U1112 ( .A(n904), .B(n110), .Z(n1248) );
  BFSVTX2 U1113 ( .A(n1886), .Z(n132) );
  EO3SVTX8 U1114 ( .A(n827), .B(n828), .C(n80), .Z(n1580) );
  NR2SVTX4 U1115 ( .A(n699), .B(n571), .Z(n1850) );
  ND2SVTX4 U1116 ( .A(n1803), .B(n1804), .Z(n1411) );
  NR2SVTX4 U1117 ( .A(n1600), .B(n1634), .Z(n1804) );
  BFSVTX12 U1118 ( .A(n1628), .Z(n497) );
  IVSVTX10 U1119 ( .A(n795), .Z(n933) );
  BFSVTX6 U1120 ( .A(m1[21]), .Z(n1060) );
  NR2SVTX4 U1121 ( .A(n233), .B(n242), .Z(n237) );
  BFSVTX1 U1122 ( .A(n414), .Z(n134) );
  EN3SVTX8 U1123 ( .A(n904), .B(n957), .C(n916), .Z(n1071) );
  NR2SVTX6 U1124 ( .A(n360), .B(n552), .Z(n185) );
  ND2SVTX4 U1125 ( .A(n139), .B(n391), .Z(n350) );
  AO6SVTX8 U1126 ( .A(n73), .B(n913), .C(n912), .Z(n307) );
  ND2SVTX4 U1127 ( .A(n515), .B(n1258), .Z(n364) );
  IVSVTX10 U1128 ( .A(n593), .Z(n838) );
  IVSVTX4 U1129 ( .A(n1982), .Z(n866) );
  IVSVTX4 U1130 ( .A(n1315), .Z(n392) );
  ND2ASVTX8 U1131 ( .A(n274), .B(n919), .Z(n1315) );
  IVSVTX6 U1132 ( .A(n950), .Z(n475) );
  ND2SVTX4 U1133 ( .A(n904), .B(n121), .Z(n152) );
  MUX21SVTX4 U1134 ( .A(n513), .B(n1137), .S(n285), .Z(n173) );
  IVSVTX12 U1135 ( .A(n869), .Z(n716) );
  ENSVTX8 U1136 ( .A(n752), .B(n1029), .Z(n1030) );
  ND4SVTX8 U1137 ( .A(n1314), .B(n2032), .C(n2030), .D(n742), .Z(n1250) );
  ND2ASVTX8 U1138 ( .A(n144), .B(n1135), .Z(n1498) );
  IVSVTX4 U1139 ( .A(n1134), .Z(n144) );
  ND3ASVTX8 U1140 ( .A(n62), .B(n231), .C(n594), .Z(n238) );
  AO20SVTX8 U1141 ( .A(n1843), .B(n753), .C(n1841), .D(n1886), .Z(n857) );
  NR2SVTX4 U1142 ( .A(m1[20]), .B(n566), .Z(n316) );
  BFSVTX6 U1143 ( .A(n909), .Z(n145) );
  NR2SVTX4 U1144 ( .A(n71), .B(n679), .Z(n1506) );
  ND3SVTX8 U1145 ( .A(n848), .B(n1516), .C(n729), .Z(n1513) );
  AO6CSVTX8 U1146 ( .A(n360), .B(n1547), .C(n1561), .Z(n1565) );
  AO7SVTX8 U1147 ( .A(n1592), .B(m1[6]), .C(n497), .Z(n662) );
  EN3SVTX8 U1148 ( .A(m1[14]), .B(m1[16]), .C(n19), .Z(n1352) );
  ND2ASVTX8 U1149 ( .A(n960), .B(n649), .Z(n653) );
  AO7SVTX4 U1150 ( .A(n704), .B(n588), .C(n116), .Z(n586) );
  EO3SVTX8 U1151 ( .A(n701), .B(n963), .C(n859), .Z(n1432) );
  ND2SVTX4 U1152 ( .A(n104), .B(n109), .Z(n864) );
  NR2SVTX4 U1153 ( .A(n917), .B(n317), .Z(n1255) );
  IVSVTX6 U1154 ( .A(n828), .Z(n735) );
  ND2SVTX4 U1155 ( .A(n1359), .B(n147), .Z(n474) );
  ND2SVTX4 U1156 ( .A(n1360), .B(n1358), .Z(n147) );
  BFSVTX1 U1157 ( .A(n535), .Z(n148) );
  BFSVTX1 U1158 ( .A(n1799), .Z(n149) );
  ND2SVTX4 U1159 ( .A(n306), .B(n1214), .Z(n1958) );
  AO6SVTX6 U1160 ( .A(n1297), .B(n1296), .C(n281), .Z(n1298) );
  AO7SVTX8 U1161 ( .A(n1637), .B(n1634), .C(n1635), .Z(n1805) );
  IVSVTX6 U1162 ( .A(n1250), .Z(n1207) );
  ND2SVTX4 U1163 ( .A(n809), .B(n1174), .Z(n309) );
  AO3ABSVTX6 U1164 ( .A(n50), .B(n265), .C(n935), .D(n544), .Z(n304) );
  ND3ABSVTX8 U1165 ( .A(n1171), .B(n282), .C(n729), .Z(n698) );
  AO7SVTX4 U1166 ( .A(n785), .B(n2), .C(n736), .Z(n778) );
  AO6SVTX6 U1167 ( .A(n1912), .B(n767), .C(n1342), .Z(n1998) );
  AO7SVTX8 U1168 ( .A(n1459), .B(n925), .C(n924), .Z(n1394) );
  NR2SVTX4 U1169 ( .A(n391), .B(n139), .Z(n351) );
  BFSVTX10 U1170 ( .A(n776), .Z(n153) );
  AO7SVTX4 U1171 ( .A(n2017), .B(n817), .C(n2012), .Z(n268) );
  IVSVTX4 U1172 ( .A(n1779), .Z(n433) );
  AO3ASVTX6 U1173 ( .A(n675), .B(n579), .C(n192), .D(n573), .Z(n213) );
  AO3CSVTX6 U1174 ( .A(n1678), .B(n1685), .C(n1865), .D(n157), .Z(n820) );
  ND3SVTX2 U1175 ( .A(n1489), .B(n717), .C(n106), .Z(n609) );
  NR2ASVTX6 U1176 ( .A(m1[23]), .B(n600), .Z(n1112) );
  NR2SVTX4 U1177 ( .A(n991), .B(n158), .Z(n992) );
  ND2SVTX4 U1178 ( .A(n159), .B(n989), .Z(n158) );
  IVSVTX4 U1179 ( .A(n990), .Z(n159) );
  AO6SVTX8 U1180 ( .A(n1979), .B(n1978), .C(n160), .Z(n1475) );
  AO7SVTX8 U1181 ( .A(n79), .B(n1531), .C(n1047), .Z(n219) );
  F_ENSVTX2 U1182 ( .A(n163), .B(n1521), .Z(n1522) );
  NR2SVTX4 U1183 ( .A(m1[0]), .B(n895), .Z(n1843) );
  AO7SVTX2 U1184 ( .A(n2029), .B(n1631), .C(n1630), .Z(n1632) );
  ND3ABSVTX8 U1185 ( .A(n851), .B(n1411), .C(n1412), .Z(n1153) );
  ND2SVTX6 U1186 ( .A(n1061), .B(n1062), .Z(n176) );
  ND3SVTX4 U1187 ( .A(n1516), .B(n117), .C(n729), .Z(n674) );
  BFSVTX1 U1188 ( .A(n1811), .Z(n166) );
  AO7ABSVTX4 U1189 ( .A(n507), .B(n526), .C(n116), .Z(n948) );
  ND2SVTX4 U1190 ( .A(n145), .B(n904), .Z(n325) );
  NR2SVTX4 U1191 ( .A(n1523), .B(n1484), .Z(n1485) );
  ND2SVTX4 U1192 ( .A(n916), .B(n669), .Z(n1005) );
  ND2ASVTX8 U1193 ( .A(n167), .B(n497), .Z(n1635) );
  IVSVTX6 U1194 ( .A(n277), .Z(n491) );
  AO17ASVTX8 U1195 ( .A(n292), .B(n287), .C(n288), .D(n1146), .Z(n1181) );
  IVSVTX4 U1196 ( .A(n816), .Z(n1656) );
  AO7SVTX2 U1197 ( .A(n790), .B(n1009), .C(n741), .Z(n1478) );
  AO3SVTX6 U1198 ( .A(n1452), .B(n380), .C(n379), .D(n63), .Z(n1418) );
  AO7SVTX8 U1199 ( .A(n863), .B(n1447), .C(n170), .Z(n1412) );
  EO3SVTX8 U1200 ( .A(n657), .B(n527), .C(n966), .Z(n1663) );
  ND3ASVTX8 U1201 ( .A(n470), .B(n182), .C(n882), .Z(n1241) );
  IVSVTX4 U1202 ( .A(n1241), .Z(n463) );
  IVSVTX4 U1203 ( .A(n783), .Z(n172) );
  BFSVTX2 U1204 ( .A(n1974), .Z(n197) );
  F_ENSVTX2 U1205 ( .A(n759), .B(n439), .Z(n438) );
  IVSVTX8 U1206 ( .A(n199), .Z(n362) );
  IVSVTX8 U1207 ( .A(n698), .Z(n806) );
  ND4ABSVTX8 U1208 ( .A(n173), .B(n698), .C(n283), .D(n1138), .Z(n1139) );
  AO6CSVTX8 U1209 ( .A(n563), .B(n929), .C(n441), .Z(n1272) );
  IVSVTX4 U1210 ( .A(n340), .Z(n736) );
  ND2SVTX4 U1211 ( .A(n933), .B(n668), .Z(n340) );
  AO7SVTX8 U1212 ( .A(n574), .B(n577), .C(n806), .Z(n192) );
  AO5NSVTX8 U1213 ( .A(n947), .B(n1592), .C(n143), .Z(n1224) );
  IVSVTX4 U1214 ( .A(n1224), .Z(n942) );
  IVSVTX10 U1215 ( .A(m1[8]), .Z(n705) );
  ND2SVTX6 U1216 ( .A(n673), .B(n687), .Z(n686) );
  ND2SVTX6 U1217 ( .A(n906), .B(n1207), .Z(n908) );
  IVSVTX4 U1218 ( .A(n177), .Z(n797) );
  EN3SVTX8 U1219 ( .A(n1140), .B(n695), .C(n145), .Z(n798) );
  IVSVTX4 U1220 ( .A(n894), .Z(n1895) );
  AO3SVTX4 U1221 ( .A(n128), .B(n1835), .C(n1834), .D(n1833), .Z(m2[9]) );
  AO7SVTX2 U1222 ( .A(n1814), .B(n1813), .C(n725), .Z(n1815) );
  ND2SVTX4 U1223 ( .A(n565), .B(n471), .Z(n182) );
  IVSVTX4 U1224 ( .A(n1540), .Z(n1551) );
  AO7SVTX6 U1225 ( .A(n1850), .B(n1849), .C(n1852), .Z(n1688) );
  ND2SVTX4 U1226 ( .A(n1572), .B(n187), .Z(n186) );
  IVSVTX4 U1227 ( .A(n205), .Z(n187) );
  IVSVTX6 U1228 ( .A(n853), .Z(n571) );
  AO7ABSVTX4 U1229 ( .A(n635), .B(n1236), .C(n1233), .Z(n1234) );
  AO7SVTX8 U1230 ( .A(n483), .B(n482), .C(n1945), .Z(n461) );
  ND4ABSVTX8 U1231 ( .A(n786), .B(n784), .C(n107), .D(n315), .Z(n805) );
  ND2ASVTX8 U1232 ( .A(n340), .B(n805), .Z(n847) );
  AO7ABSVTX4 U1233 ( .A(n1308), .B(n1651), .C(n190), .Z(n1311) );
  BFSVTX12 U1234 ( .A(n537), .Z(n265) );
  ND2SVTX8 U1235 ( .A(n96), .B(n987), .Z(n466) );
  NR2SVTX6 U1236 ( .A(n797), .B(n796), .Z(n1068) );
  IVSVTX6 U1237 ( .A(n1265), .Z(n611) );
  EOSVTX8 U1238 ( .A(n717), .B(n546), .Z(n301) );
  NR2SVTX4 U1239 ( .A(m1[6]), .B(n963), .Z(n1744) );
  NR2SVTX4 U1240 ( .A(n1578), .B(n1434), .Z(n643) );
  AO7SVTX6 U1241 ( .A(n194), .B(n193), .C(n1227), .Z(n1239) );
  IVSVTX4 U1242 ( .A(n651), .Z(n194) );
  AO7ABSVTX6 U1243 ( .A(n686), .B(n1646), .C(n1970), .Z(n1274) );
  ND2ASVTX8 U1244 ( .A(n195), .B(n945), .Z(n1222) );
  AO7SVTX6 U1245 ( .A(n335), .B(n943), .C(n1622), .Z(n195) );
  ND2SVTX4 U1246 ( .A(m1[3]), .B(m1[0]), .Z(n968) );
  ND2SVTX4 U1247 ( .A(n895), .B(m1[5]), .Z(n896) );
  IVSVTX6 U1248 ( .A(m1[20]), .Z(n807) );
  EN3SVTX8 U1249 ( .A(m1[13]), .B(n897), .C(n143), .Z(n945) );
  ND3SVTX4 U1250 ( .A(n674), .B(n1597), .C(n1513), .Z(n1196) );
  IVSVTX6 U1251 ( .A(n1185), .Z(n1302) );
  AO17SVTX8 U1252 ( .A(n1152), .B(n1153), .C(n364), .D(n363), .Z(n199) );
  BFSVTX8 U1253 ( .A(n1183), .Z(n287) );
  ND3ABSVTX8 U1254 ( .A(n1084), .B(n794), .C(n1183), .Z(n994) );
  ND3SVTX8 U1255 ( .A(n1180), .B(n217), .C(n1179), .Z(n1193) );
  ND3SVTX8 U1256 ( .A(n1136), .B(n1137), .C(n265), .Z(n1138) );
  IVSVTX4 U1257 ( .A(n238), .Z(n234) );
  IVSVTX6 U1258 ( .A(n1183), .Z(n1483) );
  ENSVTX8 U1259 ( .A(n201), .B(n1655), .Z(m2[21]) );
  NR2SVTX2 U1260 ( .A(n1650), .B(n1651), .Z(n201) );
  ND2SVTX4 U1261 ( .A(n202), .B(n1562), .Z(n1536) );
  AO7SVTX8 U1262 ( .A(n592), .B(n322), .C(n325), .Z(n799) );
  ENSVTX8 U1263 ( .A(n581), .B(n580), .Z(n687) );
  IVSVTX6 U1264 ( .A(m1[5]), .Z(n776) );
  IVSVTX2 U1265 ( .A(n1027), .Z(n206) );
  AO6SVTX2 U1266 ( .A(n1952), .B(n1953), .C(n208), .Z(n440) );
  ND2SVTX4 U1267 ( .A(n860), .B(n384), .Z(n1759) );
  ND3SVTX8 U1268 ( .A(n1118), .B(n401), .C(n399), .Z(n327) );
  AO3CDSVTX8 U1269 ( .A(n611), .B(n1268), .C(n618), .D(n698), .Z(n610) );
  AO6SVTX6 U1270 ( .A(n1257), .B(n515), .C(n514), .Z(n363) );
  ND2ASVTX8 U1271 ( .A(n1264), .B(n1498), .Z(n1265) );
  NR2SVTX4 U1272 ( .A(n400), .B(n213), .Z(n399) );
  AO6SVTX6 U1273 ( .A(n74), .B(n1147), .C(n1124), .Z(n1125) );
  NR2SVTX4 U1274 ( .A(n701), .B(n813), .Z(n1609) );
  AO6SVTX6 U1275 ( .A(n635), .B(n1236), .C(n1235), .Z(n1238) );
  IVSVTX4 U1276 ( .A(n951), .Z(n216) );
  EN3SVTX8 U1277 ( .A(m1[13]), .B(n813), .C(m1[14]), .Z(n951) );
  ND2SVTX4 U1278 ( .A(n1488), .B(n1160), .Z(n217) );
  ND3ABSVTX8 U1279 ( .A(n727), .B(n320), .C(n318), .Z(n619) );
  ND3SVTX8 U1280 ( .A(n462), .B(n530), .C(n1119), .Z(n675) );
  F_ND2ASVTX2 U1281 ( .A(n112), .B(n1162), .Z(n1163) );
  F_ENSVTX2 U1282 ( .A(n1101), .B(n219), .Z(n386) );
  NR2SVTX4 U1283 ( .A(n916), .B(n592), .Z(n1129) );
  ND2ASVTX8 U1284 ( .A(n1506), .B(n369), .Z(n1548) );
  ND2SVTX4 U1285 ( .A(n1549), .B(n1548), .Z(n1550) );
  AO7SVTX6 U1286 ( .A(n1856), .B(n1859), .C(n1857), .Z(n1694) );
  NR2SVTX4 U1287 ( .A(m1[0]), .B(n657), .Z(n1859) );
  ND2SVTX4 U1288 ( .A(n221), .B(n232), .Z(n1180) );
  F_ENSVTX2 U1289 ( .A(n74), .B(n1149), .Z(n221) );
  ND2SVTX4 U1290 ( .A(n841), .B(n426), .Z(n224) );
  AO6CSVTX8 U1291 ( .A(n73), .B(n1000), .C(n1557), .Z(n329) );
  IVSVTX8 U1292 ( .A(n572), .Z(n917) );
  ND3SVTX8 U1293 ( .A(n1577), .B(n1575), .C(n1576), .Z(m2[25]) );
  NR3SVTX8 U1294 ( .A(n1550), .B(n1563), .C(n1508), .Z(n1572) );
  IVSVTX4 U1295 ( .A(n240), .Z(n236) );
  IVSVTX12 U1296 ( .A(n321), .Z(n1488) );
  ND2SVTX6 U1297 ( .A(n933), .B(n883), .Z(n787) );
  ND2SVTX4 U1298 ( .A(n543), .B(n1481), .Z(n249) );
  F_ENSVTX2 U1299 ( .A(n763), .B(n328), .Z(n252) );
  ND2SVTX4 U1300 ( .A(n258), .B(n557), .Z(n257) );
  ND2SVTX4 U1301 ( .A(n556), .B(n1279), .Z(n258) );
  ND2SVTX4 U1302 ( .A(n89), .B(n941), .Z(n1392) );
  NR2SVTX4 U1303 ( .A(n507), .B(n77), .Z(n1395) );
  ND2SVTX4 U1304 ( .A(n1819), .B(n1391), .Z(n927) );
  ND2SVTX4 U1305 ( .A(n920), .B(n77), .Z(n1819) );
  IVSVTX4 U1306 ( .A(n713), .Z(n711) );
  ND2SVTX4 U1307 ( .A(n1612), .B(n712), .Z(n260) );
  AO20SVTX8 U1308 ( .A(n410), .B(n130), .C(n409), .D(n1129), .Z(n262) );
  AO7SVTX8 U1309 ( .A(n410), .B(n411), .C(n409), .Z(n412) );
  ND2SVTX6 U1310 ( .A(n263), .B(n264), .Z(n1130) );
  ND2SVTX6 U1311 ( .A(n1329), .B(n267), .Z(n272) );
  CTIVSVTX4 U1312 ( .A(n537), .Z(n1527) );
  ND3SVTX8 U1313 ( .A(n271), .B(n272), .C(n1134), .Z(n537) );
  ND2SVTX6 U1314 ( .A(n1462), .B(n269), .Z(n271) );
  NR2SVTX8 U1315 ( .A(n268), .B(n273), .Z(n1134) );
  ND2SVTX4 U1316 ( .A(n272), .B(n271), .Z(n270) );
  ND2ASVTX8 U1317 ( .A(n821), .B(n820), .Z(n1462) );
  IVSVTX4 U1318 ( .A(n270), .Z(n1135) );
  AO20SVTX8 U1319 ( .A(n2013), .B(n2021), .C(n1370), .D(n824), .Z(n273) );
  ND2ASVTX8 U1320 ( .A(m1[16]), .B(n473), .Z(n333) );
  ND2ASVTX8 U1321 ( .A(n897), .B(n473), .Z(n1326) );
  CTIVSVTX4 U1322 ( .A(n275), .Z(n344) );
  AO7SVTX8 U1323 ( .A(n394), .B(n2034), .C(n343), .Z(n275) );
  AO6SVTX8 U1324 ( .A(n275), .B(n906), .C(n905), .Z(n907) );
  CTBUFSVTX2 U1325 ( .A(n1462), .Z(n276) );
  ND2ASVTX8 U1326 ( .A(n950), .B(n121), .Z(n2031) );
  IVSVTX4 U1327 ( .A(n278), .Z(n1351) );
  AO5SVTX4 U1328 ( .A(n491), .B(n683), .C(n475), .Z(n278) );
  ND2ASVTX8 U1329 ( .A(n588), .B(n838), .Z(n535) );
  NR2SVTX4 U1330 ( .A(n910), .B(n340), .Z(n280) );
  ND2ASVTX8 U1331 ( .A(n1518), .B(n847), .Z(n729) );
  ND4SVTX4 U1332 ( .A(n509), .B(n1135), .C(n284), .D(n1134), .Z(n283) );
  ND2SVTX6 U1333 ( .A(n337), .B(n958), .Z(n1215) );
  AO7ABSVTX8 U1334 ( .A(n522), .B(n494), .C(n627), .Z(n1183) );
  IVSVTX8 U1335 ( .A(n523), .Z(n627) );
  ND3SVTX8 U1336 ( .A(n755), .B(n1341), .C(n652), .Z(n494) );
  AO21SVTX8 U1337 ( .A(n1244), .B(n291), .C(n1183), .D(n289), .Z(n288) );
  AO20SVTX4 U1338 ( .A(n1531), .B(n1532), .C(n1533), .D(n1597), .Z(n293) );
  ND2ASVTX8 U1339 ( .A(n593), .B(n114), .Z(n1263) );
  ND2SVTX2 U1340 ( .A(m1[16]), .B(n869), .Z(n1251) );
  ND3ASVTX6 U1341 ( .A(n1140), .B(n838), .C(n429), .Z(n428) );
  ND4SVTX8 U1342 ( .A(n304), .B(n305), .C(n302), .D(n300), .Z(n358) );
  ND2ASVTX8 U1343 ( .A(n299), .B(n303), .Z(n302) );
  AO17ASVTX8 U1344 ( .A(n797), .B(n517), .C(n313), .D(n312), .Z(n345) );
  ND3SVTX6 U1345 ( .A(n797), .B(n554), .C(n798), .Z(n312) );
  IVSVTX4 U1346 ( .A(n796), .Z(n313) );
  ND2ASVTX8 U1347 ( .A(n799), .B(n798), .Z(n517) );
  IVSVTX4 U1348 ( .A(n785), .Z(n315) );
  ND2SVTX4 U1349 ( .A(n317), .B(n316), .Z(n784) );
  ND2SVTX4 U1350 ( .A(n843), .B(n909), .Z(n320) );
  ND2SVTX8 U1351 ( .A(n1186), .B(n1275), .Z(n987) );
  NR2SVTX8 U1352 ( .A(n1182), .B(n1068), .Z(n1275) );
  NR2ASVTX8 U1353 ( .A(n799), .B(n798), .Z(n1182) );
  ND2SVTX8 U1354 ( .A(n324), .B(n323), .Z(n1186) );
  ND2SVTX8 U1355 ( .A(n916), .B(n76), .Z(n326) );
  NR2SVTX4 U1356 ( .A(n1097), .B(n79), .Z(n1051) );
  ND2SVTX4 U1357 ( .A(n111), .B(n1046), .Z(n1052) );
  NR2SVTX4 U1358 ( .A(n916), .B(n119), .Z(n1045) );
  IVSVTX4 U1359 ( .A(n189), .Z(n387) );
  ND2ASVTX8 U1360 ( .A(n389), .B(n327), .Z(n398) );
  AO6SVTX4 U1361 ( .A(n1008), .B(n746), .C(n1007), .Z(n328) );
  ND3SVTX6 U1362 ( .A(n1102), .B(n99), .C(n181), .Z(n1095) );
  AO20SVTX8 U1363 ( .A(n332), .B(n330), .C(n1075), .D(n1074), .Z(n1102) );
  IVSVTX4 U1364 ( .A(n331), .Z(n330) );
  IVSVTX12 U1365 ( .A(n869), .Z(n1140) );
  ND2SVTX4 U1366 ( .A(n475), .B(n957), .Z(n338) );
  AN2SVTX8 U1367 ( .A(n278), .B(n339), .Z(n628) );
  IVSVTX12 U1368 ( .A(m1[17]), .Z(n572) );
  ND2ASVTX8 U1369 ( .A(n1199), .B(n1201), .Z(n1167) );
  CTIVSVTX4 U1370 ( .A(n559), .Z(n511) );
  IVSVTX8 U1371 ( .A(m1[21]), .Z(n909) );
  AO1CSVTX6 U1372 ( .A(n994), .B(n992), .C(n94), .D(n939), .Z(n346) );
  IVSVTX4 U1373 ( .A(n350), .Z(n1856) );
  NR2SVTX6 U1374 ( .A(n352), .B(n1836), .Z(n1886) );
  IVSVTX4 U1375 ( .A(n351), .Z(n1857) );
  ND2SVTX4 U1376 ( .A(n1836), .B(n352), .Z(n1885) );
  ND2ASVTX8 U1377 ( .A(n352), .B(m1[6]), .Z(n825) );
  ND2ASVTX8 U1378 ( .A(n1092), .B(n536), .Z(n567) );
  NR2SVTX8 U1379 ( .A(n1546), .B(n1545), .Z(m2[24]) );
  ND2SVTX8 U1380 ( .A(n708), .B(n1191), .Z(n402) );
  NR2SVTX8 U1381 ( .A(n1552), .B(n1569), .Z(n1539) );
  IVSVTX8 U1382 ( .A(n1547), .Z(n1569) );
  NR2ASVTX6 U1383 ( .A(n1535), .B(n354), .Z(n1552) );
  ND2ASVTX8 U1384 ( .A(n1535), .B(n354), .Z(n1547) );
  IVSVTX12 U1385 ( .A(m1[14]), .Z(n473) );
  ND3ABSVTX8 U1386 ( .A(m1[27]), .B(m1[26]), .C(n356), .Z(n1171) );
  NR2SVTX8 U1387 ( .A(n1510), .B(n1651), .Z(n626) );
  NR3ABSVTX6 U1388 ( .A(n1306), .B(n624), .C(n357), .Z(n1651) );
  ND2SVTX8 U1389 ( .A(n1549), .B(n1548), .Z(n1553) );
  IVSVTX12 U1390 ( .A(n362), .Z(n1008) );
  AO6SVTX8 U1391 ( .A(n508), .B(n1115), .C(n370), .Z(n1557) );
  ND2SVTX4 U1392 ( .A(n990), .B(n76), .Z(n1114) );
  AO7SVTX6 U1393 ( .A(n1148), .B(n1120), .C(n1122), .Z(n1115) );
  NR2SVTX4 U1394 ( .A(n1112), .B(n1022), .Z(n508) );
  NR2SVTX4 U1395 ( .A(n910), .B(n916), .Z(n1022) );
  NR3SVTX8 U1396 ( .A(n695), .B(n91), .C(n88), .Z(n892) );
  ND2ASVTX8 U1397 ( .A(n777), .B(n116), .Z(n1918) );
  IVSVTX4 U1398 ( .A(n1323), .Z(n371) );
  F_ENSVTX2 U1399 ( .A(n1372), .B(n373), .Z(n372) );
  AO7SVTX6 U1400 ( .A(n381), .B(n1713), .C(n376), .Z(n1454) );
  ND2SVTX4 U1401 ( .A(n860), .B(n32), .Z(n376) );
  AO6ASVTX8 U1402 ( .A(n383), .B(n1418), .C(n377), .Z(n604) );
  ND2SVTX4 U1403 ( .A(n607), .B(n1454), .Z(n379) );
  ND2ASVTX8 U1404 ( .A(n1628), .B(n384), .Z(n1747) );
  AO7ABSVTX8 U1405 ( .A(n117), .B(n1516), .C(n385), .Z(n1597) );
  ND2SVTX4 U1406 ( .A(n543), .B(n386), .Z(n464) );
  ND2SVTX4 U1407 ( .A(n1978), .B(n212), .Z(n1980) );
  NR2SVTX4 U1408 ( .A(n391), .B(m1[6]), .Z(n816) );
  NR2SVTX6 U1409 ( .A(n1093), .B(n536), .Z(n444) );
  NR2SVTX8 U1410 ( .A(n396), .B(n395), .Z(n1541) );
  NR2SVTX8 U1411 ( .A(n397), .B(n444), .Z(n1653) );
  ND2ASVTX8 U1412 ( .A(n81), .B(n583), .Z(n1118) );
  MUX21NSVTX8 U1413 ( .A(n591), .B(n590), .S(n582), .Z(n401) );
  ND3SVTX8 U1414 ( .A(n415), .B(n417), .C(n416), .Z(n1191) );
  IVSVTX4 U1415 ( .A(n507), .Z(n405) );
  NR2SVTX6 U1416 ( .A(n950), .B(n584), .Z(n1906) );
  ND2SVTX4 U1417 ( .A(n588), .B(n592), .Z(n2003) );
  IVSVTX4 U1418 ( .A(n2005), .Z(n407) );
  ND2ASVTX8 U1419 ( .A(n572), .B(n116), .Z(n2005) );
  AO6CSVTX8 U1420 ( .A(n1906), .B(n1337), .C(n1336), .Z(n1365) );
  ND2SVTX4 U1421 ( .A(n2002), .B(n2004), .Z(n930) );
  ND2SVTX4 U1422 ( .A(n457), .B(m1[3]), .Z(n1896) );
  ND2SVTX8 U1423 ( .A(n419), .B(n418), .Z(n1573) );
  ND3SVTX8 U1424 ( .A(n1973), .B(n1969), .C(n1274), .Z(n418) );
  NR2SVTX6 U1425 ( .A(n1974), .B(n1644), .Z(n419) );
  ND2SVTX6 U1426 ( .A(n422), .B(n1573), .Z(n1654) );
  ND2SVTX4 U1427 ( .A(n1612), .B(n1614), .Z(n1821) );
  ND2SVTX4 U1428 ( .A(n777), .B(n963), .Z(n1612) );
  ND2SVTX4 U1429 ( .A(n841), .B(n432), .Z(n425) );
  NR2SVTX4 U1430 ( .A(n1060), .B(n76), .Z(n486) );
  NR2SVTX4 U1431 ( .A(n430), .B(n428), .Z(n709) );
  ND2ASVTX8 U1432 ( .A(n431), .B(n919), .Z(n430) );
  NR2ASVTX6 U1433 ( .A(n473), .B(n839), .Z(n432) );
  NR2ASVTX6 U1434 ( .A(n433), .B(n455), .Z(n841) );
  ND2SVTX4 U1435 ( .A(n181), .B(n542), .Z(n991) );
  AO17SVTX4 U1436 ( .A(n1253), .B(n102), .C(n437), .D(n1254), .Z(n436) );
  AO7SVTX6 U1437 ( .A(n1252), .B(n344), .C(n1251), .Z(n437) );
  NR3SVTX8 U1438 ( .A(m1[0]), .B(n1836), .C(n842), .Z(n844) );
  ND2SVTX4 U1439 ( .A(n445), .B(n31), .Z(n842) );
  IVSVTX4 U1440 ( .A(n837), .Z(n448) );
  NR2SVTX4 U1441 ( .A(n86), .B(n847), .Z(n449) );
  ENSVTX8 U1442 ( .A(n1131), .B(n1130), .Z(n451) );
  ND3SVTX6 U1443 ( .A(n458), .B(n454), .C(n453), .Z(n694) );
  NR2SVTX4 U1444 ( .A(n842), .B(n839), .Z(n453) );
  ND2SVTX8 U1445 ( .A(n456), .B(n457), .Z(n455) );
  IVSVTX8 U1446 ( .A(m1[6]), .Z(n457) );
  NR4SVTX8 U1447 ( .A(n630), .B(n571), .C(m1[0]), .D(n89), .Z(n458) );
  IVSVTX4 U1448 ( .A(n839), .Z(n840) );
  ND2SVTX4 U1449 ( .A(n699), .B(n496), .Z(n1713) );
  ND2SVTX6 U1450 ( .A(n735), .B(n496), .Z(n734) );
  ND2SVTX4 U1451 ( .A(n564), .B(n461), .Z(n1970) );
  NR2ASVTX4 U1452 ( .A(n1273), .B(n461), .Z(n1243) );
  AO7ABSVTX4 U1453 ( .A(n708), .B(n1191), .C(n398), .Z(n1508) );
  ND2SVTX6 U1454 ( .A(n1284), .B(n1424), .Z(n1094) );
  ND4SVTX4 U1455 ( .A(n841), .B(n840), .C(n844), .D(n468), .Z(n471) );
  IVSVTX4 U1456 ( .A(n920), .Z(n683) );
  IVSVTX4 U1457 ( .A(n474), .Z(n1984) );
  ND2SVTX4 U1458 ( .A(n473), .B(m1[16]), .Z(n1358) );
  ND2SVTX4 U1459 ( .A(m1[14]), .B(n919), .Z(n1359) );
  ENSVTX4 U1460 ( .A(n1082), .B(n1081), .Z(n583) );
  AO6SVTX8 U1461 ( .A(n1008), .B(n1042), .C(n1041), .Z(n1043) );
  ND4ABSVTX8 U1462 ( .A(n76), .B(n699), .C(n479), .D(n476), .Z(n540) );
  NR3SVTX6 U1463 ( .A(m1[16]), .B(n478), .C(n477), .Z(n476) );
  IVSVTX12 U1464 ( .A(m1[15]), .Z(n950) );
  AO7SVTX8 U1465 ( .A(n1239), .B(n1238), .C(n100), .Z(n1962) );
  ND2SVTX6 U1466 ( .A(n1234), .B(n650), .Z(n1961) );
  ND2ASVTX8 U1467 ( .A(n560), .B(n481), .Z(n1945) );
  AO6SVTX8 U1468 ( .A(n1961), .B(n1962), .C(n914), .Z(n482) );
  ND2SVTX4 U1469 ( .A(n70), .B(n484), .Z(n1273) );
  NR2SVTX4 U1470 ( .A(n733), .B(n1196), .Z(n484) );
  CTIVSVTX4 U1471 ( .A(n910), .Z(n485) );
  ND4SVTX4 U1472 ( .A(n487), .B(n511), .C(n105), .D(n892), .Z(n489) );
  NR2SVTX4 U1473 ( .A(n1077), .B(n1094), .Z(n490) );
  IVSVTX4 U1474 ( .A(n232), .Z(n1424) );
  ND2SVTX4 U1475 ( .A(n277), .B(n1140), .Z(n1249) );
  ND2SVTX4 U1476 ( .A(n89), .B(n491), .Z(n956) );
  AO7SVTX6 U1477 ( .A(n89), .B(n491), .C(n917), .Z(n955) );
  ND2ASVTX8 U1478 ( .A(n822), .B(n1826), .Z(n1325) );
  AN2SVTX8 U1479 ( .A(n1620), .B(n743), .Z(n1826) );
  ND2SVTX4 U1480 ( .A(n522), .B(n494), .Z(n521) );
  IVSVTX4 U1481 ( .A(n495), .Z(n750) );
  ND2SVTX8 U1482 ( .A(n496), .B(n77), .Z(n500) );
  ND2SVTX4 U1483 ( .A(n1010), .B(n412), .Z(n550) );
  ND2SVTX4 U1484 ( .A(n897), .B(n80), .Z(n1824) );
  ND2SVTX4 U1485 ( .A(n80), .B(n630), .Z(n1768) );
  ND2SVTX4 U1486 ( .A(n508), .B(n1116), .Z(n1517) );
  IVSVTX4 U1487 ( .A(n509), .Z(n1137) );
  ND2SVTX2 U1488 ( .A(m1[16]), .B(n918), .Z(n1210) );
  AO7SVTX8 U1489 ( .A(n868), .B(n1984), .C(n867), .Z(n1257) );
  ND2SVTX4 U1490 ( .A(n518), .B(n1075), .Z(n1187) );
  NR2SVTX8 U1491 ( .A(n964), .B(n1578), .Z(n984) );
  NR2SVTX8 U1492 ( .A(n519), .B(n979), .Z(n1578) );
  ND2SVTX8 U1493 ( .A(n663), .B(n662), .Z(n731) );
  EO3SVTX8 U1494 ( .A(m1[11]), .B(n677), .C(n1592), .Z(n979) );
  ND2SVTX8 U1495 ( .A(n521), .B(n627), .Z(n580) );
  NR2SVTX8 U1496 ( .A(n1228), .B(n985), .Z(n522) );
  AO7SVTX8 U1497 ( .A(n1998), .B(n985), .C(n524), .Z(n523) );
  IVSVTX4 U1498 ( .A(n813), .Z(n525) );
  AN2SVTX8 U1499 ( .A(m1[11]), .B(n162), .Z(n1634) );
  IVSVTX12 U1500 ( .A(m1[7]), .Z(n827) );
  ND2SVTX4 U1501 ( .A(n630), .B(n493), .Z(n1743) );
  NR2SVTX4 U1502 ( .A(m1[7]), .B(n1830), .Z(n1741) );
  IVSVTX4 U1503 ( .A(n695), .Z(n601) );
  NR2SVTX4 U1504 ( .A(n669), .B(n1501), .Z(n1556) );
  ND2SVTX4 U1505 ( .A(n933), .B(n911), .Z(n1501) );
  NR2SVTX4 U1506 ( .A(n701), .B(n77), .Z(n1600) );
  ND2SVTX4 U1507 ( .A(n1937), .B(n849), .Z(n851) );
  ND2SVTX4 U1508 ( .A(n953), .B(n954), .Z(n1910) );
  ND2SVTX4 U1509 ( .A(n952), .B(n951), .Z(n1386) );
  NR2SVTX8 U1510 ( .A(n1909), .B(n533), .Z(n767) );
  NR2SVTX8 U1511 ( .A(n953), .B(n954), .Z(n1909) );
  NR2SVTX6 U1512 ( .A(n944), .B(n945), .Z(n531) );
  ND4SVTX8 U1513 ( .A(n1066), .B(n1067), .C(n1065), .D(n1064), .Z(n536) );
  ND3ABSVTX6 U1514 ( .A(n1104), .B(n1492), .C(n537), .Z(n538) );
  NR2SVTX8 U1515 ( .A(n669), .B(n281), .Z(n544) );
  ND2SVTX4 U1516 ( .A(n548), .B(n547), .Z(n1195) );
  ND2SVTX4 U1517 ( .A(n88), .B(n1140), .Z(n551) );
  ND2SVTX6 U1518 ( .A(n93), .B(n1571), .Z(n552) );
  ND2SVTX8 U1519 ( .A(n1562), .B(n553), .Z(n1571) );
  ND2SVTX8 U1520 ( .A(n568), .B(n567), .Z(n1563) );
  NR2SVTX4 U1521 ( .A(m1[27]), .B(m1[26]), .Z(n889) );
  NR2ASVTX6 U1522 ( .A(n1952), .B(n672), .Z(n932) );
  NR2SVTX4 U1523 ( .A(m1[6]), .B(n860), .Z(n722) );
  IVSVTX2 U1524 ( .A(m1[6]), .Z(n859) );
  ND2SVTX8 U1525 ( .A(n562), .B(n1992), .Z(n985) );
  NR2SVTX8 U1526 ( .A(n656), .B(n1217), .Z(n562) );
  NR2ASVTX8 U1527 ( .A(n655), .B(n958), .Z(n1217) );
  AO7SVTX6 U1528 ( .A(n1353), .B(n628), .C(n1350), .Z(n1995) );
  ND2SVTX4 U1529 ( .A(n118), .B(n586), .Z(n960) );
  ND2SVTX4 U1530 ( .A(n473), .B(n593), .Z(n2032) );
  EO3SVTX8 U1531 ( .A(n566), .B(n588), .C(n592), .Z(n1218) );
  ND2SVTX4 U1532 ( .A(m1[14]), .B(n572), .Z(n2033) );
  ND2SVTX6 U1533 ( .A(n576), .B(n575), .Z(n574) );
  ND3ABSVTX8 U1534 ( .A(n1182), .B(n1185), .C(n1183), .Z(n582) );
  IVSVTX4 U1535 ( .A(n897), .Z(n584) );
  ND2SVTX4 U1536 ( .A(n588), .B(n585), .Z(n1324) );
  IVSVTX4 U1537 ( .A(n920), .Z(n585) );
  ND2SVTX4 U1538 ( .A(n950), .B(n918), .Z(n2002) );
  ND2SVTX4 U1539 ( .A(n910), .B(n1526), .Z(n596) );
  NR2SVTX4 U1540 ( .A(n1140), .B(n601), .Z(n1120) );
  ND2SVTX4 U1541 ( .A(n695), .B(n807), .Z(n599) );
  ND2SVTX4 U1542 ( .A(n601), .B(n600), .Z(n1079) );
  IVSVTX4 U1543 ( .A(n807), .Z(n600) );
  ND2SVTX4 U1544 ( .A(n601), .B(n136), .Z(n1122) );
  ND4SVTX4 U1545 ( .A(n990), .B(n601), .C(n1529), .D(n781), .Z(n1197) );
  NR2SVTX4 U1546 ( .A(n355), .B(n941), .Z(n898) );
  NR3SVTX8 U1547 ( .A(n92), .B(n1563), .C(n608), .Z(n1509) );
  NR2SVTX4 U1548 ( .A(n1267), .B(n1265), .Z(n612) );
  IVSVTX4 U1549 ( .A(n616), .Z(n613) );
  ND2SVTX4 U1550 ( .A(n1488), .B(n1261), .Z(n614) );
  ND2SVTX2 U1551 ( .A(n917), .B(n728), .Z(n617) );
  EO3SVTX8 U1552 ( .A(n950), .B(n897), .C(n355), .Z(n954) );
  AO7SVTX6 U1553 ( .A(n622), .B(n621), .C(n620), .Z(n1177) );
  NR2SVTX4 U1554 ( .A(n670), .B(n1527), .Z(n622) );
  IVSVTX4 U1555 ( .A(n625), .Z(n623) );
  ND2SVTX4 U1556 ( .A(n1188), .B(n1483), .Z(n1189) );
  NR2SVTX4 U1557 ( .A(n140), .B(n630), .Z(n1658) );
  IVSVTX4 U1558 ( .A(n629), .Z(n1464) );
  ND2SVTX4 U1559 ( .A(n630), .B(n966), .Z(n629) );
  ND2SVTX4 U1560 ( .A(n106), .B(n660), .Z(n631) );
  IVSVTX4 U1561 ( .A(n660), .Z(n632) );
  NR2SVTX4 U1562 ( .A(n803), .B(n633), .Z(n660) );
  ND3SVTX6 U1563 ( .A(n635), .B(n122), .C(n1341), .Z(n1994) );
  ND4ABSVTX8 U1564 ( .A(n637), .B(n975), .C(n1581), .D(n636), .Z(n652) );
  IVSVTX4 U1565 ( .A(n654), .Z(n636) );
  NR2SVTX4 U1566 ( .A(n1441), .B(n967), .Z(n1581) );
  NR2SVTX4 U1567 ( .A(n1437), .B(n691), .Z(n637) );
  F_ENSVTX2 U1568 ( .A(n2001), .B(n642), .Z(n641) );
  AO7SVTX6 U1569 ( .A(n648), .B(n1434), .C(n1662), .Z(n1440) );
  NR2SVTX8 U1570 ( .A(n978), .B(n977), .Z(n1434) );
  ND2SVTX8 U1571 ( .A(n978), .B(n977), .Z(n1662) );
  IVSVTX4 U1572 ( .A(n1441), .Z(n645) );
  NR2SVTX4 U1573 ( .A(n967), .B(n964), .Z(n646) );
  ND2SVTX6 U1574 ( .A(n1664), .B(n1663), .Z(n648) );
  IVSVTX4 U1575 ( .A(n961), .Z(n649) );
  NR2SVTX8 U1576 ( .A(n100), .B(n1239), .Z(n650) );
  ND2SVTX4 U1577 ( .A(n651), .B(n1993), .Z(n1235) );
  NR3SVTX8 U1578 ( .A(n561), .B(n1989), .C(n628), .Z(n651) );
  ND2SVTX6 U1579 ( .A(n1915), .B(n767), .Z(n1228) );
  NR2SVTX4 U1580 ( .A(m1[1]), .B(n657), .Z(n753) );
  ND2SVTX4 U1581 ( .A(n232), .B(n1522), .Z(n659) );
  ND2SVTX8 U1582 ( .A(n800), .B(n64), .Z(n1072) );
  ND2SVTX6 U1583 ( .A(n984), .B(n1582), .Z(n661) );
  ND2SVTX4 U1584 ( .A(n408), .B(n1592), .Z(n663) );
  IVSVTX4 U1585 ( .A(n849), .Z(n664) );
  ND2SVTX4 U1586 ( .A(m1[25]), .B(m1[26]), .Z(n893) );
  NR2SVTX4 U1587 ( .A(n1033), .B(n1104), .Z(n1287) );
  NR2ASVTX6 U1588 ( .A(n791), .B(n916), .Z(n1033) );
  F_ENSVTX2 U1589 ( .A(n1008), .B(n1132), .Z(n1141) );
  BFSVTX12 U1590 ( .A(m1[5]), .Z(n966) );
  IVSVTX8 U1591 ( .A(n791), .Z(n668) );
  IVSVTX10 U1592 ( .A(n915), .Z(n669) );
  AO7SVTX2 U1593 ( .A(n1283), .B(n1282), .C(n1281), .Z(n1306) );
  F_ND2ASVTX2 U1594 ( .A(m1[10]), .B(n827), .Z(n692) );
  AO6SVTX2 U1595 ( .A(n2009), .B(n1954), .C(n1953), .Z(n1955) );
  ND2SVTX4 U1596 ( .A(n1167), .B(n937), .Z(n1240) );
  AO7SVTX1 U1597 ( .A(n722), .B(n726), .C(n24), .Z(n1760) );
  AN2ABSVTX4 U1598 ( .A(n1217), .B(n1216), .Z(n1237) );
  F_ND2SVTX1 U1599 ( .A(n2031), .B(n2030), .Z(n2039) );
  AO1ABSVTX4 U1600 ( .A(n1208), .B(n1207), .C(n1206), .D(n1205), .Z(n1209) );
  NR2SVTX4 U1601 ( .A(n1507), .B(n1551), .Z(n1512) );
  ND2ASVTX8 U1602 ( .A(n97), .B(n681), .Z(n680) );
  NR2SVTX4 U1603 ( .A(n699), .B(n496), .Z(n682) );
  IVSVTX4 U1604 ( .A(n1089), .Z(n1085) );
  AO7CSVTX4 U1605 ( .A(n1502), .B(n1557), .C(n1556), .Z(n1503) );
  AO7SVTX6 U1606 ( .A(n1648), .B(n1971), .C(n1647), .Z(n1977) );
  NR2SVTX0H U1607 ( .A(n722), .B(n1757), .Z(n1761) );
  NR2ASVTX6 U1608 ( .A(n391), .B(n433), .Z(n684) );
  ND2SVTX4 U1609 ( .A(n701), .B(n966), .Z(n1721) );
  IVSVTX2 U1610 ( .A(n1412), .Z(n688) );
  IVSVTX2 U1611 ( .A(n686), .Z(n690) );
  NR2SVTX0H U1612 ( .A(n1264), .B(n1946), .Z(n1947) );
  F_IVSVTX0H U1613 ( .A(n59), .Z(n1772) );
  IVSVTX2 U1614 ( .A(n1517), .Z(n1000) );
  IVSVTX12 U1615 ( .A(m1[20]), .Z(n904) );
  IVSVTX2 U1616 ( .A(n1235), .Z(n1233) );
  ND2SVTX2 U1617 ( .A(n1337), .B(n1336), .Z(n1339) );
  ND2SVTX4 U1618 ( .A(n806), .B(n1038), .Z(n1066) );
  ND2SVTX2 U1619 ( .A(n1962), .B(n1961), .Z(n1963) );
  ND2SVTX4 U1620 ( .A(n699), .B(n527), .Z(n1706) );
  NR2SVTX2 U1621 ( .A(n1102), .B(n1096), .Z(n1077) );
  ND3SVTX4 U1622 ( .A(n819), .B(n1846), .C(n972), .Z(n976) );
  ND2SVTX2 U1623 ( .A(n1303), .B(n580), .Z(n1304) );
  ND2SVTX4 U1624 ( .A(n1907), .B(n1337), .Z(n700) );
  ND2SVTX4 U1625 ( .A(n393), .B(n777), .Z(n1907) );
  FAS1SVTX4 U1626 ( .A(n668), .B(n933), .CI(n76), .CO(n802), .Z(n796) );
  AO3ABSVTX6 U1627 ( .A(n707), .B(n1531), .C(n1058), .D(n1057), .Z(n1063) );
  ND2SVTX4 U1628 ( .A(n145), .B(n136), .Z(n744) );
  AN2ABSVTX6 U1629 ( .A(n909), .B(n12), .Z(n1123) );
  ND2SVTX4 U1630 ( .A(m1[26]), .B(n915), .Z(n887) );
  AO6SVTX2 U1631 ( .A(n1259), .B(n1258), .C(n1257), .Z(n1260) );
  ND2SVTX4 U1632 ( .A(n467), .B(n1482), .Z(n1301) );
  FAS1SVTX4 U1633 ( .A(n916), .B(n119), .CI(n915), .CO(n792), .Z(n793) );
  ND2SVTX2 U1634 ( .A(n909), .B(n12), .Z(n1148) );
  ND3ABSVTX1 U1635 ( .A(n1171), .B(n1174), .C(n1170), .Z(n1176) );
  OR2SVTX4 U1636 ( .A(n918), .B(m1[16]), .Z(n749) );
  ENSVTX4 U1637 ( .A(n1972), .B(n1971), .Z(m2[16]) );
  ENSVTX4 U1638 ( .A(n1977), .B(n1976), .Z(m2[17]) );
  IVSVTX2 U1639 ( .A(n732), .Z(n733) );
  ND2ASVTX8 U1640 ( .A(n1569), .B(n1570), .Z(n1564) );
  NR3SVTX2 U1641 ( .A(n1250), .B(n1203), .C(n604), .Z(n1206) );
  AN2SVTX4 U1642 ( .A(n895), .B(n776), .Z(n739) );
  IVSVTX2 U1643 ( .A(n1068), .Z(n1070) );
  NR2SVTX2 U1644 ( .A(n998), .B(n1517), .Z(n913) );
  ND2SVTX2 U1645 ( .A(n696), .B(n772), .Z(n1867) );
  ND2SVTX4 U1646 ( .A(n1152), .B(n1153), .Z(n1259) );
  ND2SVTX2 U1647 ( .A(n1796), .B(n1225), .Z(n1226) );
  ND2SVTX4 U1648 ( .A(n1783), .B(n826), .Z(n1327) );
  IVSVTX2 U1649 ( .A(n1990), .Z(n1220) );
  AO6CSVTX2 U1650 ( .A(n1008), .B(n57), .C(n744), .Z(n1081) );
  AO7SVTX6 U1651 ( .A(n1078), .B(n744), .C(n1079), .Z(n1041) );
  IVSVTX4 U1652 ( .A(n1496), .Z(n1109) );
  IVSVTX2 U1653 ( .A(n808), .Z(n811) );
  AO7SVTX2 U1654 ( .A(n1494), .B(n1493), .C(n11), .Z(n1495) );
  IVSVTX4 U1655 ( .A(m1[26]), .Z(n837) );
  NR2SVTX2 U1656 ( .A(n569), .B(n1983), .Z(n1212) );
  IVSVTX2 U1657 ( .A(n1059), .Z(n707) );
  F_ND2SVTX0H U1658 ( .A(n47), .B(n629), .Z(n1729) );
  IVSVTX2 U1659 ( .A(n563), .Z(n1820) );
  ND3SVTX1 U1660 ( .A(n2016), .B(n2015), .C(n2014), .Z(n2020) );
  IVSVTX2 U1661 ( .A(n1051), .Z(n1054) );
  IVSVTX2 U1662 ( .A(n1524), .Z(n873) );
  IVSVTX2 U1663 ( .A(n1527), .Z(n1297) );
  AO7SVTX2 U1664 ( .A(n1295), .B(n1293), .C(n1288), .Z(n1292) );
  IVSVTX6 U1665 ( .A(n1531), .Z(n1056) );
  NR2SVTX2 U1666 ( .A(n129), .B(n1530), .Z(n1533) );
  ND2SVTX2 U1667 ( .A(n225), .B(n1592), .Z(n1593) );
  F_ENSVTX2 U1668 ( .A(n756), .B(n1213), .Z(n1214) );
  IVSVTX2 U1669 ( .A(n580), .Z(n1282) );
  AO6SVTX2 U1670 ( .A(n1482), .B(n345), .C(n1277), .Z(n1278) );
  B_ND2SVTX1 U1671 ( .A(m1[0]), .B(n203), .Z(n1838) );
  F_EOSVTX2 U1672 ( .A(n1456), .B(n1455), .Z(n1457) );
  AO7SVTX2 U1673 ( .A(n1737), .B(n1585), .C(n45), .Z(n1586) );
  B_ND2SVTX2 U1674 ( .A(n1392), .B(n1391), .Z(n1399) );
  ND2SVTX2 U1675 ( .A(n543), .B(n1369), .Z(n1374) );
  ND2SVTX2 U1676 ( .A(n1088), .B(n1089), .Z(n1090) );
  ND2SVTX4 U1677 ( .A(n1086), .B(n1085), .Z(n1091) );
  F_EOSVTX2 U1678 ( .A(n1988), .B(n1987), .Z(n2042) );
  B_ND2SVTX0H U1679 ( .A(n1970), .B(n1969), .Z(n1972) );
  IVSVTX2 U1680 ( .A(n1572), .Z(n1567) );
  AO6ABSVTX8 U1681 ( .A(n1568), .B(n1567), .C(n1566), .Z(m2[26]) );
  AO6SVTX2 U1682 ( .A(n1599), .B(n1718), .C(n1598), .Z(n1605) );
  NR2SVTX2 U1683 ( .A(n1106), .B(n1492), .Z(n1107) );
  NR3SVTX2 U1684 ( .A(n1087), .B(n466), .C(n82), .Z(n1088) );
  AO6SVTX8 U1685 ( .A(n1099), .B(n84), .C(n934), .Z(n1009) );
  NR2ASVTX6 U1686 ( .A(n91), .B(n807), .Z(n810) );
  AO7ABSVTX2 U1687 ( .A(n543), .B(n2027), .C(n2026), .Z(n2028) );
  ND3SVTX4 U1688 ( .A(n1302), .B(n1184), .C(n1183), .Z(n1190) );
  AO4SVTX2 U1689 ( .A(n1538), .B(n1537), .C(n1551), .D(n1539), .Z(n1544) );
  NR2ASVTX6 U1690 ( .A(n1309), .B(n1312), .Z(n1310) );
  ND2SVTX2 U1691 ( .A(n1060), .B(n1240), .Z(n1061) );
  ND2SVTX2 U1692 ( .A(n1140), .B(n917), .Z(n800) );
  IVSVTX2 U1693 ( .A(n942), .Z(n962) );
  AO1SVTX8 U1694 ( .A(n1313), .B(n1312), .C(n1311), .D(n1310), .Z(m2[22]) );
  IVSVTX2 U1695 ( .A(n889), .Z(n1013) );
  ND2SVTX2 U1696 ( .A(n917), .B(n76), .Z(n1270) );
  NR2SVTX2 U1697 ( .A(m1[24]), .B(m1[27]), .Z(n781) );
  ND3SVTX4 U1698 ( .A(n1092), .B(n1091), .C(n1090), .Z(n1093) );
  F_AO2SVTX1 U1699 ( .A(n806), .B(n1839), .C(n165), .D(m1[1]), .Z(n1864) );
  AO6SVTX1 U1700 ( .A(n2025), .B(n806), .C(n762), .Z(n2026) );
  AO6SVTX1 U1701 ( .A(n1629), .B(n806), .C(n764), .Z(n1630) );
  ND3SVTX2 U1702 ( .A(n88), .B(n1200), .C(n1201), .Z(n1202) );
  F_ND2SVTX0H U1703 ( .A(n88), .B(m1[26]), .Z(n1198) );
  F_ENSVTX2 U1704 ( .A(n751), .B(n1260), .Z(n1261) );
  NR2SVTX2 U1705 ( .A(n1009), .B(n910), .Z(n1530) );
  IVSVTX2 U1706 ( .A(n1272), .Z(n2009) );
  NR2SVTX2 U1707 ( .A(n1651), .B(n1308), .Z(n1309) );
  ND2SVTX4 U1708 ( .A(n776), .B(n1779), .Z(n720) );
  AO7SVTX2 U1709 ( .A(n1255), .B(n1155), .C(n1256), .Z(n1156) );
  EOSVTX2 U1710 ( .A(n915), .B(n1060), .Z(n1489) );
  ND3ASVTX6 U1711 ( .A(n721), .B(n1541), .C(n1542), .Z(n1543) );
  F_ND2ASVTX2 U1712 ( .A(m1[7]), .B(n353), .Z(n1726) );
  EOSVTX2 U1713 ( .A(n1589), .B(n1813), .Z(n1599) );
  NR2SVTX2 U1714 ( .A(n1014), .B(n1013), .Z(n1015) );
  F_ND3SVTX2 U1715 ( .A(n1960), .B(n1959), .C(n1958), .Z(n1965) );
  IVSVTX0H U1716 ( .A(n1758), .Z(n726) );
  ND2SVTX2 U1717 ( .A(m1[0]), .B(n772), .Z(n1849) );
  B_ND2SVTX2 U1718 ( .A(n129), .B(n1627), .Z(n1534) );
  F_AO2SVTX1 U1719 ( .A(n806), .B(n1680), .C(n165), .D(n203), .Z(n1700) );
  F_AO2SVTX1 U1720 ( .A(n1718), .B(n1672), .C(n165), .D(n140), .Z(n1673) );
  AO7SVTX8 U1721 ( .A(n908), .B(n604), .C(n907), .Z(n1505) );
  AO6SVTX4 U1722 ( .A(n1259), .B(n1212), .C(n1211), .Z(n1213) );
  NR2SVTX2 U1723 ( .A(m1[0]), .B(m1[3]), .Z(n969) );
  IVSVTX4 U1724 ( .A(n1288), .Z(n730) );
  IVSVTX2 U1725 ( .A(n1493), .Z(n1288) );
  ND2SVTX2 U1726 ( .A(n988), .B(n466), .Z(n989) );
  NR2SVTX2 U1727 ( .A(m1[26]), .B(m1[27]), .Z(n1017) );
  NR2SVTX2 U1728 ( .A(n1252), .B(n1250), .Z(n1253) );
  ND2SVTX2 U1729 ( .A(n742), .B(n1314), .Z(n1378) );
  OR2SVTX6 U1730 ( .A(n704), .B(n393), .Z(n742) );
  OR2ABSVTX4 U1731 ( .A(m1[20]), .B(m1[23]), .Z(n1098) );
  IVSVTX4 U1732 ( .A(n737), .Z(n738) );
  ND3SVTX4 U1733 ( .A(n1560), .B(n1012), .C(n81), .Z(n1561) );
  ND2SVTX2 U1734 ( .A(n1836), .B(n699), .Z(n1868) );
  ND2SVTX2 U1735 ( .A(m1[1]), .B(n699), .Z(n1852) );
  NR2SVTX2 U1736 ( .A(n699), .B(n527), .Z(n1668) );
  ND2SVTX4 U1737 ( .A(n777), .B(n1830), .Z(n1404) );
  IVSVTX4 U1738 ( .A(n819), .Z(n1685) );
  ND2SVTX2 U1739 ( .A(n772), .B(n696), .Z(n974) );
  NR2SVTX2 U1740 ( .A(n1556), .B(n1518), .Z(n1519) );
  NR2SVTX2 U1741 ( .A(n1039), .B(n1004), .Z(n746) );
  IVSVTX2 U1742 ( .A(n1167), .Z(n1168) );
  ND2ASVTX8 U1743 ( .A(n919), .B(n592), .Z(n1266) );
  ND2SVTX2 U1744 ( .A(n566), .B(n1140), .Z(n1262) );
  FAS1SVTX4 U1745 ( .A(n716), .B(m1[16]), .CI(n957), .CO(n940), .Z(n958) );
  ND2SVTX4 U1746 ( .A(n1302), .B(n1275), .Z(n1084) );
  FAS1SVTX4 U1747 ( .A(m1[6]), .B(n391), .CI(n1779), .CO(n981), .Z(n977) );
  ND2SVTX2 U1748 ( .A(n232), .B(n740), .Z(n1560) );
  FAS1SVTX4 U1749 ( .A(n699), .B(n1836), .CI(n966), .CO(n1664), .Z(n1437) );
  ND2SVTX4 U1750 ( .A(n1549), .B(n997), .Z(n1308) );
  IVSVTX8 U1751 ( .A(n915), .Z(n990) );
  AO6SVTX4 U1752 ( .A(n1542), .B(n1541), .C(n1536), .Z(n1546) );
  ND2SVTX2 U1753 ( .A(n1547), .B(n1573), .Z(n1568) );
  ND2SVTX4 U1754 ( .A(n1361), .B(n21), .Z(n1983) );
  NR2SVTX2 U1755 ( .A(n695), .B(n910), .Z(n1001) );
  BFSVTX12 U1756 ( .A(m1[21]), .Z(n916) );
  OR2SVTX4 U1757 ( .A(n1197), .B(n837), .Z(n937) );
  F_ND2SVTX0H U1758 ( .A(n911), .B(n1554), .Z(n1555) );
  ND2SVTX2 U1759 ( .A(n695), .B(n910), .Z(n1003) );
  AO4SVTX2 U1760 ( .A(n1050), .B(n1048), .C(n1049), .D(n1052), .Z(n1058) );
  IVSVTX4 U1761 ( .A(n1099), .Z(n1047) );
  ND2SVTX2 U1762 ( .A(n736), .B(n786), .Z(n780) );
  IVSVTX8 U1763 ( .A(n706), .Z(n860) );
  ND2ASVTX8 U1764 ( .A(n1204), .B(n344), .Z(n1208) );
  BFSVTX12 U1765 ( .A(m1[12]), .Z(n897) );
  AO6NSVTX1 U1766 ( .A(n1504), .B(n74), .C(n1558), .Z(n740) );
  ENSVTX0H U1767 ( .A(n1318), .B(n1317), .Z(n747) );
  ENSVTX0H U1768 ( .A(n1590), .B(n1820), .Z(n748) );
  AN2SVTX0H U1769 ( .A(n1210), .B(n749), .Z(n756) );
  AO7SVTX6 U1770 ( .A(n1127), .B(n1161), .C(n1128), .Z(n1099) );
  AN2SVTX0H U1771 ( .A(n910), .B(m1[26]), .Z(n757) );
  F_ND2ASVTX2 U1772 ( .A(n1140), .B(n916), .Z(n1080) );
  AN2SVTX0H U1773 ( .A(n123), .B(n1627), .Z(n764) );
  OR2SVTX1 U1774 ( .A(n1198), .B(n1197), .Z(n765) );
  AN2SVTX0H U1775 ( .A(m1[11]), .B(n1627), .Z(n770) );
  NR2SVTX2 U1776 ( .A(n353), .B(m1[3]), .Z(n1883) );
  IVSVTX2 U1777 ( .A(n1883), .Z(n856) );
  AO7SVTX4 U1778 ( .A(n876), .B(n875), .C(n874), .Z(n877) );
  AN2BSVTX4 U1779 ( .A(n1484), .B(n876), .Z(n872) );
  IVSVTX4 U1780 ( .A(n1523), .Z(n876) );
  IVSVTX4 U1781 ( .A(n107), .Z(n775) );
  IVSVTX12 U1782 ( .A(n895), .Z(n1836) );
  NR2SVTX4 U1783 ( .A(n933), .B(n792), .Z(n804) );
  IVSVTX4 U1784 ( .A(n812), .Z(n1370) );
  ND2SVTX4 U1785 ( .A(n735), .B(n525), .Z(n1622) );
  IVSVTX4 U1786 ( .A(n814), .Z(n1403) );
  ND2SVTX4 U1787 ( .A(n963), .B(n526), .Z(n1620) );
  ND2SVTX4 U1788 ( .A(n1656), .B(n1726), .Z(n1463) );
  ND2SVTX4 U1789 ( .A(n860), .B(n527), .Z(n1783) );
  AO7SVTX2 U1790 ( .A(n1868), .B(n1865), .C(n1867), .Z(n821) );
  NR2SVTX2 U1791 ( .A(m1[1]), .B(n772), .Z(n818) );
  NR3ABSVTX2 U1792 ( .A(m1[0]), .B(n1836), .C(n818), .Z(n1678) );
  ND2SVTX2 U1793 ( .A(n701), .B(m1[6]), .Z(n1784) );
  ND2SVTX4 U1794 ( .A(n630), .B(n497), .Z(n1780) );
  NR2SVTX6 U1795 ( .A(n669), .B(n1060), .Z(n1039) );
  NR2SVTX4 U1796 ( .A(n1039), .B(n1001), .Z(n871) );
  ND2SVTX4 U1797 ( .A(n599), .B(n1080), .Z(n1004) );
  IVSVTX4 U1798 ( .A(n1004), .Z(n1042) );
  ND2SVTX4 U1799 ( .A(n871), .B(n1042), .Z(n1524) );
  ND2SVTX4 U1800 ( .A(n701), .B(n493), .Z(n1637) );
  NR2SVTX6 U1801 ( .A(n722), .B(n1754), .Z(n862) );
  NR2SVTX4 U1802 ( .A(n1704), .B(n1668), .Z(n1756) );
  ND2SVTX4 U1803 ( .A(n1756), .B(n862), .Z(n863) );
  AO20SVTX8 U1804 ( .A(n858), .B(n857), .C(n856), .D(n855), .Z(n1447) );
  ND2SVTX4 U1805 ( .A(n963), .B(n630), .Z(n1755) );
  NR2SVTX4 U1806 ( .A(n904), .B(n957), .Z(n1150) );
  NR2ASVTX6 U1807 ( .A(n1484), .B(n873), .Z(n875) );
  ND3SVTX2 U1808 ( .A(m1[26]), .B(m1[25]), .C(n890), .Z(n886) );
  ND2SVTX4 U1809 ( .A(n701), .B(n526), .Z(n1608) );
  ND2SVTX2 U1810 ( .A(n897), .B(n950), .Z(n1929) );
  NR2SVTX4 U1811 ( .A(n1123), .B(n1120), .Z(n1116) );
  NR2SVTX4 U1812 ( .A(n1140), .B(n695), .Z(n1127) );
  NR2SVTX8 U1813 ( .A(n700), .B(n930), .Z(n1954) );
  ND2ASVTX8 U1814 ( .A(n947), .B(n209), .Z(n1614) );
  NR2SVTX4 U1815 ( .A(n1821), .B(n927), .Z(n929) );
  ND2SVTX2 U1816 ( .A(m1[3]), .B(m1[6]), .Z(n1875) );
  ND2SVTX4 U1817 ( .A(n957), .B(n916), .Z(n1161) );
  AO7SVTX4 U1818 ( .A(n1098), .B(n1045), .C(n1046), .Z(n934) );
  IVSVTX4 U1819 ( .A(n813), .Z(n941) );
  EN3SVTX8 U1820 ( .A(n963), .B(n941), .C(n704), .Z(n1223) );
  ND2ASVTX8 U1821 ( .A(n942), .B(n1223), .Z(n1797) );
  ND2SVTX4 U1822 ( .A(n949), .B(n948), .Z(n953) );
  ND2SVTX4 U1823 ( .A(n956), .B(n955), .Z(n1219) );
  ND2SVTX6 U1824 ( .A(n1219), .B(n1218), .Z(n1990) );
  ND2SVTX4 U1825 ( .A(n1351), .B(n1352), .Z(n1350) );
  FAS1SVTX4 U1826 ( .A(m1[5]), .B(n701), .CI(n1779), .CO(n1433), .Z(n1442) );
  IVSVTX4 U1827 ( .A(n1848), .Z(n971) );
  AO7SVTX2 U1828 ( .A(n772), .B(n696), .C(m1[6]), .Z(n973) );
  ND2SVTX4 U1829 ( .A(n974), .B(n973), .Z(n978) );
  ND2SVTX4 U1830 ( .A(n731), .B(n1580), .Z(n1738) );
  ND2SVTX4 U1831 ( .A(n980), .B(n979), .Z(n1579) );
  IVSVTX4 U1832 ( .A(n1442), .Z(n982) );
  IVSVTX0H U1833 ( .A(n998), .Z(n999) );
  IVSVTX0H U1834 ( .A(n1001), .Z(n1002) );
  IVSVTX0H U1835 ( .A(n1022), .Z(n1024) );
  NR2SVTX2 U1836 ( .A(n1112), .B(n1025), .Z(n1028) );
  AO7SVTX2 U1837 ( .A(n1112), .B(n1026), .C(n1114), .Z(n1027) );
  ND2ASVTX8 U1838 ( .A(n299), .B(n1030), .Z(n1067) );
  IVSVTX0H U1839 ( .A(n1039), .Z(n1040) );
  ND2SVTX4 U1840 ( .A(n1056), .B(n1055), .Z(n1057) );
  ND2ASVTX8 U1841 ( .A(n1084), .B(n580), .Z(n1089) );
  NR2SVTX4 U1842 ( .A(n1105), .B(n1104), .Z(n1106) );
  IVSVTX0H U1843 ( .A(n1112), .Z(n1113) );
  IVSVTX0H U1844 ( .A(n1120), .Z(n1121) );
  ND2SVTX4 U1845 ( .A(n1143), .B(n101), .Z(n1145) );
  NR2SVTX2 U1846 ( .A(n1255), .B(n1154), .Z(n1157) );
  IVSVTX2 U1847 ( .A(n1257), .Z(n1155) );
  IVSVTX2 U1848 ( .A(n1215), .Z(n1216) );
  ND3SVTX2 U1849 ( .A(n1224), .B(n1223), .C(n1222), .Z(n1225) );
  IVSVTX4 U1850 ( .A(n1440), .Z(n1230) );
  NR2SVTX4 U1851 ( .A(n1231), .B(n1232), .Z(n1236) );
  IVSVTX4 U1852 ( .A(n1243), .Z(n1969) );
  IVSVTX0H U1853 ( .A(n1246), .Z(n1247) );
  ND2SVTX2 U1854 ( .A(n1248), .B(n1247), .Z(n1254) );
  IVSVTX0H U1855 ( .A(n672), .Z(n1269) );
  ND2SVTX8 U1856 ( .A(n421), .B(n1654), .Z(n1312) );
  NR2SVTX2 U1857 ( .A(n1295), .B(n1289), .Z(n1290) );
  AO7SVTX2 U1858 ( .A(n420), .B(n1651), .C(n169), .Z(n1307) );
  ND2SVTX2 U1859 ( .A(n1314), .B(n1315), .Z(n1318) );
  ENSVTX0H U1860 ( .A(n1321), .B(n1320), .Z(n1335) );
  AO7SVTX1 U1861 ( .A(n188), .B(n1920), .C(n1918), .Z(n1330) );
  AO8SVTX1 U1862 ( .A(n2016), .B(n1326), .C(n2015), .D(n1330), .Z(n1331) );
  ENSVTX0H U1863 ( .A(n1332), .B(n1331), .Z(n1333) );
  AO6SVTX1 U1864 ( .A(n2009), .B(n1907), .C(n1906), .Z(n1338) );
  EOSVTX0H U1865 ( .A(n1339), .B(n1338), .Z(n1347) );
  IVSVTX0H U1866 ( .A(n561), .Z(n1355) );
  AO6SVTX1 U1867 ( .A(n1994), .B(n676), .C(n1912), .Z(n1343) );
  AO7SVTX2 U1868 ( .A(n142), .B(n1343), .C(n737), .Z(n1344) );
  F_ENSVTX2 U1869 ( .A(n1345), .B(n1344), .Z(n1346) );
  AO2SVTX2 U1870 ( .A(n1347), .B(n543), .C(n673), .D(n1346), .Z(n1348) );
  AO7SVTX1 U1871 ( .A(n1352), .B(n1351), .C(n1350), .Z(n1357) );
  AO7SVTX1 U1872 ( .A(n1998), .B(n561), .C(n18), .Z(n1354) );
  AO6SVTX1 U1873 ( .A(n1320), .B(n1361), .C(n1360), .Z(n1362) );
  EOSVTX2 U1874 ( .A(n1363), .B(n1362), .Z(n1364) );
  NR2ASVTX1 U1875 ( .A(n2017), .B(n2018), .Z(n1372) );
  ND2SVTX4 U1876 ( .A(n1385), .B(n1384), .Z(m2[13]) );
  NR2ASVTX1 U1877 ( .A(n1386), .B(n533), .Z(n1389) );
  IVSVTX0H U1878 ( .A(n1821), .Z(n1393) );
  AO6SVTX1 U1879 ( .A(n1819), .B(n713), .C(n1395), .Z(n1396) );
  AO7SVTX1 U1880 ( .A(n1397), .B(n1820), .C(n1396), .Z(n1398) );
  ENSVTX0H U1881 ( .A(n1399), .B(n1398), .Z(n1400) );
  NR2SVTX1 U1882 ( .A(n1403), .B(n1402), .Z(n1409) );
  IVSVTX0H U1883 ( .A(n1404), .Z(n1405) );
  AO7SVTX1 U1884 ( .A(n1406), .B(n1405), .C(n1824), .Z(n1407) );
  AO8SVTX1 U1885 ( .A(n1826), .B(n689), .C(n2015), .D(n1407), .Z(n1408) );
  ENSVTX0H U1886 ( .A(n1409), .B(n1408), .Z(n1410) );
  AO6SVTX1 U1887 ( .A(n1410), .B(n806), .C(n770), .Z(n1428) );
  BFSVTX1 U1888 ( .A(n1411), .Z(n1932) );
  BFSVTX1 U1889 ( .A(n1413), .Z(n1934) );
  AO7SVTX1 U1890 ( .A(n1932), .B(n688), .C(n1934), .Z(n1414) );
  ENSVTX0H U1891 ( .A(n1415), .B(n1414), .Z(n1426) );
  IVSVTX0H U1892 ( .A(n1418), .Z(n1813) );
  AO6SVTX1 U1893 ( .A(n1419), .B(n166), .C(n902), .Z(n1420) );
  AO7SVTX1 U1894 ( .A(n1432), .B(n1433), .C(n1431), .Z(n1445) );
  IVSVTX0H U1895 ( .A(n1846), .Z(n1439) );
  NR2SVTX2 U1896 ( .A(n1439), .B(n1438), .Z(n1687) );
  ND2SVTX2 U1897 ( .A(n1685), .B(n52), .Z(n1684) );
  AO17ASVTX4 U1898 ( .A(n52), .B(n819), .C(n1687), .D(n1684), .Z(n1892) );
  AO8ASVTX4 U1899 ( .A(n60), .B(n1890), .C(n1892), .D(n1440), .Z(n1701) );
  AO7SVTX2 U1900 ( .A(n1701), .B(n7), .C(n1443), .Z(n1444) );
  ND2SVTX2 U1901 ( .A(n852), .B(n24), .Z(n1449) );
  IVSVTX0H U1902 ( .A(n1447), .Z(n1762) );
  AO6SVTX1 U1903 ( .A(n1762), .B(n23), .C(n1758), .Z(n1448) );
  EOSVTX0H U1904 ( .A(n1449), .B(n1448), .Z(n1450) );
  IVSVTX0H U1905 ( .A(n1452), .Z(n1751) );
  AO6SVTX1 U1906 ( .A(n1751), .B(n1453), .C(n1746), .Z(n1455) );
  AO6SVTX1 U1907 ( .A(n1775), .B(n1769), .C(n59), .Z(n1460) );
  EOSVTX0H U1908 ( .A(n1461), .B(n1460), .Z(n1470) );
  ND2SVTX2 U1909 ( .A(n1727), .B(n47), .Z(n1465) );
  ENSVTX0H U1910 ( .A(n1467), .B(n1785), .Z(n1468) );
  AO4SVTX1 U1911 ( .A(n1322), .B(n859), .C(n1468), .D(n718), .Z(n1469) );
  ENSVTX8 U1912 ( .A(n1476), .B(n1475), .Z(m2[20]) );
  NR2SVTX2 U1913 ( .A(n790), .B(n1532), .Z(n1479) );
  NR2SVTX2 U1914 ( .A(n1523), .B(n1524), .Z(n1486) );
  ND2SVTX8 U1915 ( .A(n1573), .B(n1509), .Z(n1542) );
  AO6CSVTX8 U1916 ( .A(n1542), .B(n1541), .C(n1549), .Z(n1511) );
  ENSVTX8 U1917 ( .A(n1512), .B(n1511), .Z(m2[23]) );
  AO1ABSVTX2 U1918 ( .A(n86), .B(n1516), .C(n1515), .D(n1514), .Z(n1535) );
  NR2SVTX2 U1919 ( .A(n61), .B(n1524), .Z(n1525) );
  ND2SVTX4 U1920 ( .A(n1543), .B(n1544), .Z(n1545) );
  ND2SVTX6 U1921 ( .A(n1564), .B(n1565), .Z(n1566) );
  NR2SVTX2 U1922 ( .A(n93), .B(n1569), .Z(n1574) );
  NR2SVTX2 U1923 ( .A(n731), .B(n1580), .Z(n1737) );
  ENSVTX0H U1924 ( .A(n1591), .B(n2015), .Z(n1595) );
  AO7SVTX2 U1925 ( .A(n1597), .B(n748), .C(n1596), .Z(n1598) );
  EOSVTX0H U1926 ( .A(n1602), .B(n688), .Z(n1603) );
  AO7SVTX1 U1927 ( .A(n1609), .B(n1813), .C(n151), .Z(n1610) );
  ENSVTX0H U1928 ( .A(n1611), .B(n1610), .Z(n1643) );
  AO7SVTX1 U1929 ( .A(n1616), .B(n1820), .C(n1615), .Z(n1617) );
  ENSVTX0H U1930 ( .A(n1618), .B(n1617), .Z(n1633) );
  NR2ASVTX1 U1931 ( .A(n1797), .B(n149), .Z(n1619) );
  ENSVTX0H U1932 ( .A(n1619), .B(n1994), .Z(n1631) );
  NR2ASVTX1 U1933 ( .A(n1622), .B(n1621), .Z(n1626) );
  IVSVTX0H U1934 ( .A(n1623), .Z(n1624) );
  AO6SVTX1 U1935 ( .A(n2015), .B(n46), .C(n1624), .Z(n1625) );
  ENSVTX0H U1936 ( .A(n1626), .B(n1625), .Z(n1629) );
  ND2SVTX2 U1937 ( .A(n1636), .B(n1635), .Z(n1639) );
  AO7SVTX1 U1938 ( .A(n1600), .B(n688), .C(n1637), .Z(n1638) );
  ENSVTX0H U1939 ( .A(n1639), .B(n1638), .Z(n1640) );
  IVSVTX2 U1940 ( .A(n1969), .Z(n1648) );
  BFSVTX2 U1941 ( .A(n1970), .Z(n1647) );
  ND2SVTX2 U1942 ( .A(n825), .B(n1656), .Z(n1657) );
  ENSVTX0H U1943 ( .A(n1657), .B(n276), .Z(n1661) );
  ND2SVTX2 U1944 ( .A(n1722), .B(n1723), .Z(n1659) );
  ENSVTX0H U1945 ( .A(n1659), .B(n1775), .Z(n1660) );
  F_AO2SVTX1 U1946 ( .A(n806), .B(n1661), .C(n543), .D(n1660), .Z(n1676) );
  ENSVTX0H U1947 ( .A(n1669), .B(n1762), .Z(n1670) );
  ENSVTX0H U1948 ( .A(n1671), .B(n1751), .Z(n1672) );
  IVSVTX0H U1949 ( .A(n1868), .Z(n1677) );
  NR2SVTX2 U1950 ( .A(n1685), .B(n1678), .Z(n1869) );
  ENSVTX0H U1951 ( .A(n1679), .B(n1869), .Z(n1680) );
  EOSVTX0H U1952 ( .A(n771), .B(n1682), .Z(n1683) );
  AO7SVTX1 U1953 ( .A(n1685), .B(n52), .C(n1684), .Z(n1686) );
  IVSVTX0H U1954 ( .A(n40), .Z(n1689) );
  ND2SVTX2 U1955 ( .A(n1876), .B(n1689), .Z(n1690) );
  EOSVTX0H U1956 ( .A(n1877), .B(n1690), .Z(n1691) );
  EOSVTX0H U1957 ( .A(n1695), .B(n1897), .Z(n1696) );
  ND2SVTX2 U1958 ( .A(n1705), .B(n720), .Z(n1710) );
  AO6SVTX1 U1959 ( .A(n1762), .B(n1708), .C(n1707), .Z(n1709) );
  EOSVTX0H U1960 ( .A(n1710), .B(n1709), .Z(n1711) );
  AO6SVTX1 U1961 ( .A(n1751), .B(n1714), .C(n685), .Z(n1715) );
  AO6SVTX1 U1962 ( .A(n1775), .B(n1723), .C(n684), .Z(n1724) );
  EOSVTX0H U1963 ( .A(n1725), .B(n1724), .Z(n1732) );
  ENSVTX0H U1964 ( .A(n1729), .B(n1728), .Z(n1730) );
  AO4SVTX1 U1965 ( .A(n1322), .B(n153), .C(n1730), .D(n718), .Z(n1731) );
  IVSVTX0H U1966 ( .A(n1741), .Z(n1742) );
  ND2SVTX2 U1967 ( .A(n1743), .B(n1742), .Z(n1753) );
  IVSVTX0H U1968 ( .A(n1453), .Z(n1745) );
  IVSVTX0H U1969 ( .A(n1746), .Z(n1748) );
  AO6SVTX1 U1970 ( .A(n1751), .B(n1750), .C(n1749), .Z(n1752) );
  AO6SVTX1 U1971 ( .A(n1762), .B(n1761), .C(n1760), .Z(n1763) );
  F_AO2SVTX1 U1972 ( .A(n1766), .B(n1718), .C(n1765), .D(n678), .Z(n1793) );
  ND2SVTX2 U1973 ( .A(n1768), .B(n692), .Z(n1778) );
  IVSVTX0H U1974 ( .A(n1769), .Z(n1770) );
  IVSVTX0H U1975 ( .A(n1780), .Z(n1781) );
  F_IVSVTX1 U1976 ( .A(n1783), .Z(n1786) );
  ENSVTX0H U1977 ( .A(n1788), .B(n1787), .Z(n1789) );
  AO6SVTX2 U1978 ( .A(n543), .B(n1791), .C(n1790), .Z(n1792) );
  IVSVTX0H U1979 ( .A(n1804), .Z(n1807) );
  AO7SVTX1 U1980 ( .A(n1807), .B(n688), .C(n1806), .Z(n1808) );
  ENSVTX0H U1981 ( .A(n1809), .B(n1808), .Z(n1818) );
  AO7SVTX1 U1982 ( .A(n1821), .B(n1820), .C(n711), .Z(n1822) );
  ENSVTX0H U1983 ( .A(n1823), .B(n1822), .Z(n1832) );
  ND2SVTX2 U1984 ( .A(n1824), .B(n1404), .Z(n1828) );
  AO6SVTX1 U1985 ( .A(n2015), .B(n1826), .C(n1825), .Z(n1827) );
  ENSVTX0H U1986 ( .A(n1828), .B(n1827), .Z(n1829) );
  ENSVTX0H U1987 ( .A(n1838), .B(n1837), .Z(n1839) );
  EOSVTX0H U1988 ( .A(n1843), .B(n1842), .Z(n1844) );
  ENSVTX0H U1989 ( .A(n1848), .B(n1847), .Z(n1855) );
  IVSVTX0H U1990 ( .A(n1850), .Z(n1851) );
  EOSVTX0H U1991 ( .A(n968), .B(n1853), .Z(n1854) );
  F_AO2SVTX1 U1992 ( .A(n673), .B(n1855), .C(n543), .D(n1854), .Z(n1862) );
  ND2SVTX2 U1993 ( .A(n1857), .B(n350), .Z(n1858) );
  EOSVTX0H U1994 ( .A(n1859), .B(n1858), .Z(n1860) );
  IVSVTX0H U1995 ( .A(n1865), .Z(n1866) );
  ENSVTX0H U1996 ( .A(n1872), .B(n1871), .Z(n1882) );
  AO7SVTX1 U1997 ( .A(n40), .B(n1877), .C(n1876), .Z(n1879) );
  ENSVTX0H U1998 ( .A(n1880), .B(n1879), .Z(n1881) );
  F_AO2SVTX1 U1999 ( .A(n806), .B(n1882), .C(n543), .D(n1881), .Z(n1905) );
  ND2SVTX2 U2000 ( .A(n1884), .B(n856), .Z(n1888) );
  AO7SVTX1 U2001 ( .A(n132), .B(n771), .C(n1885), .Z(n1887) );
  ENSVTX0H U2002 ( .A(n1888), .B(n1887), .Z(n1889) );
  F_ND2ASVTX2 U2003 ( .A(n1891), .B(n1890), .Z(n1893) );
  ENSVTX0H U2004 ( .A(n1893), .B(n1892), .Z(n1894) );
  ENSVTX0H U2005 ( .A(n1900), .B(n1899), .Z(n1901) );
  ENSVTX0H U2006 ( .A(n1908), .B(n2009), .Z(n1928) );
  ND2SVTX2 U2007 ( .A(n1911), .B(n1910), .Z(n1917) );
  AO7SVTX1 U2008 ( .A(n533), .B(n1913), .C(n1386), .Z(n1914) );
  AO8SVTX2 U2009 ( .A(n1915), .B(n1994), .C(n1387), .D(n1914), .Z(n1916) );
  IVSVTX0H U2010 ( .A(n188), .Z(n1921) );
  AO6SVTX1 U2011 ( .A(n2015), .B(n2016), .C(n1921), .Z(n1922) );
  ENSVTX0H U2012 ( .A(n1923), .B(n1922), .Z(n1924) );
  ND2SVTX1 U2013 ( .A(n742), .B(n1929), .Z(n1930) );
  ENSVTX0H U2014 ( .A(n1930), .B(n102), .Z(n1943) );
  AO6SVTX1 U2015 ( .A(n1937), .B(n516), .C(n1936), .Z(n1938) );
  AO7SVTX1 U2016 ( .A(n688), .B(n1939), .C(n1938), .Z(n1940) );
  ENSVTX0H U2017 ( .A(n1941), .B(n1940), .Z(n1942) );
  F_AO2SVTX1 U2018 ( .A(n1943), .B(n1718), .C(n1942), .D(n678), .Z(n1944) );
  IVSVTX0H U2019 ( .A(n1266), .Z(n1946) );
  ENSVTX0H U2020 ( .A(n365), .B(n1947), .Z(n1951) );
  ND2SVTX2 U2021 ( .A(n543), .B(n1957), .Z(n1959) );
  NR2SVTX2 U2022 ( .A(n1965), .B(n1964), .Z(n1966) );
  ND2SVTX2 U2023 ( .A(n1982), .B(n1981), .Z(n1988) );
  IVSVTX0H U2024 ( .A(n1992), .Z(n1997) );
  IVSVTX0H U2025 ( .A(n1995), .Z(n1996) );
  AO7SVTX1 U2026 ( .A(n1998), .B(n1997), .C(n1996), .Z(n1999) );
  AO7SVTX1 U2027 ( .A(n2006), .B(n1365), .C(n2005), .Z(n2007) );
  AO6SVTX1 U2028 ( .A(n2009), .B(n2008), .C(n2007), .Z(n2010) );
  EOSVTX0H U2029 ( .A(n2011), .B(n2010), .Z(n2027) );
  ENSVTX0H U2030 ( .A(n2024), .B(n2023), .Z(n2025) );
  AO7SVTX1 U2031 ( .A(n9), .B(n2035), .C(n2033), .Z(n2036) );
  ND2SVTX2 U2032 ( .A(n1718), .B(n2040), .Z(n2041) );
endmodule


module remap_top ( num_i, rslt_o );
  input [31:0] num_i;
  output [31:0] rslt_o;
  wire   n167, n168, n169, n170, n171, n172, n174, n175, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n266, n267, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n354, n355, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n409, n410,
         n411, n412, n413, n414, n415, n416, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n513, n514, n515, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n682, n683, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750;
  wire   [27:0] keyvalues_m1;

  remap re_map ( .m1({keyvalues_m1[27:14], n465, keyvalues_m1[12:8], n468, 
        n470, keyvalues_m1[5:0]}), .m2(rslt_o[26:0]) );
  BFSVTX0H U200 ( .A(n455), .Z(rslt_o[31]) );
  AO6ASVTX4 U201 ( .A(n628), .B(n664), .C(n663), .Z(n750) );
  BFSVTX6 U202 ( .A(n312), .Z(n373) );
  AO4ABSVTX6 U203 ( .C(n327), .D(n566), .A(n648), .B(n683), .Z(n567) );
  IVSVTX10 U204 ( .A(n319), .Z(n628) );
  CTIVSVTX2 U205 ( .A(n686), .Z(n566) );
  NR4ABSVTX6 U206 ( .A(n312), .B(n742), .C(n649), .D(n743), .Z(n655) );
  CTIVSVTX2 U207 ( .A(n184), .Z(n672) );
  IVSVTX10 U208 ( .A(n438), .Z(keyvalues_m1[5]) );
  BFSVTX0H U209 ( .A(n502), .Z(n184) );
  IVSVTX10 U210 ( .A(n635), .Z(keyvalues_m1[11]) );
  ND2ASVTX6 U211 ( .A(n172), .B(n737), .Z(n330) );
  AO7SVTX1 U212 ( .A(n543), .B(n298), .C(n542), .Z(n551) );
  AO4SVTX6 U213 ( .A(n221), .B(n312), .C(n409), .D(n640), .Z(n380) );
  AO2SVTX6 U214 ( .A(n219), .B(n682), .C(n391), .D(n310), .Z(n331) );
  ND3SVTX4 U215 ( .A(n227), .B(n741), .C(n742), .Z(n744) );
  BFSVTX8 U216 ( .A(n254), .Z(n262) );
  CTBUFSVTX4 U217 ( .A(n636), .Z(n172) );
  IVSVTX0H U218 ( .A(n271), .Z(n334) );
  ND2ASVTX4 U219 ( .A(n568), .B(n683), .Z(n650) );
  AO7ASVTX6 U220 ( .A(n738), .B(n739), .C(n312), .Z(n314) );
  ND3SVTX4 U221 ( .A(n276), .B(n686), .C(n171), .Z(n647) );
  ND3ABSVTX4 U222 ( .A(n281), .B(n273), .C(n191), .Z(n690) );
  AO7SVTX2 U223 ( .A(n335), .B(rslt_o[29]), .C(n666), .Z(n670) );
  IVSVTX10 U224 ( .A(n363), .Z(n312) );
  CTBUFSVTX4 U225 ( .A(n216), .Z(n171) );
  ND2SVTX2 U226 ( .A(n454), .B(n657), .Z(n676) );
  IVSVTX0H U227 ( .A(n569), .Z(n667) );
  CTIVSVTX2 U228 ( .A(n638), .Z(n383) );
  ND2SVTX4 U229 ( .A(n572), .B(n573), .Z(n717) );
  IVSVTX0H U230 ( .A(n202), .Z(n405) );
  IVSVTX0H U231 ( .A(n689), .Z(n296) );
  ND3SVTX4 U232 ( .A(n379), .B(n484), .C(n319), .Z(n378) );
  NR2SVTX6 U233 ( .A(n277), .B(n628), .Z(n258) );
  MUX21NSVTX6 U234 ( .A(n522), .B(n728), .S(n287), .Z(n632) );
  AO2SVTX4 U235 ( .A(n644), .B(n484), .C(rslt_o[29]), .D(n390), .Z(n344) );
  AO7SVTX2 U236 ( .A(n199), .B(n709), .C(n706), .Z(n711) );
  IVSVTX2 U237 ( .A(n627), .Z(n522) );
  IVSVTX4 U238 ( .A(rslt_o[29]), .Z(n277) );
  ND2ASVTX4 U239 ( .A(n431), .B(n430), .Z(n630) );
  ND3SVTX6 U240 ( .A(n379), .B(n293), .C(n628), .Z(n210) );
  IVSVTX2 U241 ( .A(n291), .Z(n540) );
  AN2SVTX4 U242 ( .A(n230), .B(n472), .Z(n644) );
  NR2SVTX2 U243 ( .A(n492), .B(n274), .Z(n390) );
  CTIVSVTX10 U244 ( .A(n732), .Z(n253) );
  AO7SVTX4 U245 ( .A(n611), .B(n610), .C(n428), .Z(n523) );
  AO7ASVTX2 U246 ( .A(num_i[16]), .B(n475), .C(n482), .Z(n279) );
  B_ND2SVTX2 U247 ( .A(n704), .B(n637), .Z(n626) );
  NR2SVTX2 U248 ( .A(rslt_o[29]), .B(n612), .Z(n261) );
  ND3ASVTX4 U249 ( .A(n199), .B(n454), .C(n607), .Z(n423) );
  BFSVTX6 U250 ( .A(n464), .Z(n293) );
  ND3SVTX6 U251 ( .A(n600), .B(num_i[7]), .C(n274), .Z(n596) );
  NR2ASVTX2 U252 ( .A(num_i[3]), .B(n475), .Z(n488) );
  IVSVTX8 U253 ( .A(n464), .Z(n484) );
  IVSVTX4 U254 ( .A(n428), .Z(n704) );
  CTBUFSVTX4 U255 ( .A(n385), .Z(n224) );
  CTIVSVTX2 U256 ( .A(n466), .Z(n487) );
  IVSVTX0H U257 ( .A(n560), .Z(n582) );
  BFSVTX4 U258 ( .A(n389), .Z(n274) );
  CTBUFSVTX4 U259 ( .A(n472), .Z(n266) );
  NR3SVTX4 U260 ( .A(n475), .B(n202), .C(n597), .Z(n593) );
  IVSVTX6 U261 ( .A(n607), .Z(n657) );
  IVSVTX2 U262 ( .A(n591), .Z(n597) );
  IVSVTX10 U263 ( .A(n389), .Z(n475) );
  IVSVTX0H U264 ( .A(n552), .Z(n588) );
  IVSVTX2 U265 ( .A(num_i[5]), .Z(n202) );
  IVSVTX0H U266 ( .A(num_i[16]), .Z(n617) );
  IVSVTX0H U267 ( .A(n230), .Z(n594) );
  ND2ASVTX4 U268 ( .A(n668), .B(n472), .Z(n616) );
  BFSVTX2 U269 ( .A(num_i[12]), .Z(n569) );
  IVSVTX8 U270 ( .A(n267), .Z(n472) );
  IVSVTX2 U271 ( .A(num_i[8]), .Z(n668) );
  ND2ASVTX6 U272 ( .A(n485), .B(n437), .Z(n298) );
  IVSVTX6 U273 ( .A(n198), .Z(n643) );
  OR2SVTX6 U274 ( .A(n466), .B(n485), .Z(n425) );
  NR3ABSVTX6 U275 ( .A(n560), .B(n578), .C(n290), .Z(n247) );
  IVSVTX8 U276 ( .A(n364), .Z(n389) );
  IVSVTX2 U277 ( .A(n584), .Z(n578) );
  NR2ASVTX4 U278 ( .A(n192), .B(n571), .Z(n345) );
  IVSVTX8 U279 ( .A(n485), .Z(n198) );
  IVSVTX2 U280 ( .A(n514), .Z(n483) );
  IVSVTX2 U281 ( .A(n508), .Z(n471) );
  NR3SVTX6 U282 ( .A(n410), .B(n412), .C(n411), .Z(n399) );
  IVSVTX2 U283 ( .A(num_i[9]), .Z(n229) );
  CTBUFSVTX4 U284 ( .A(n538), .Z(n211) );
  BFSVTX2 U285 ( .A(num_i[10]), .Z(n586) );
  NR3SVTX4 U286 ( .A(n575), .B(n537), .C(n562), .Z(n354) );
  BFSVTX2 U287 ( .A(n469), .Z(n571) );
  OR2SVTX2 U288 ( .A(num_i[31]), .B(num_i[30]), .Z(n476) );
  ND2SVTX2 U289 ( .A(num_i[18]), .B(n495), .Z(n498) );
  CTBUFSVTX4 U290 ( .A(n194), .Z(n182) );
  CTBUFSVTX4 U291 ( .A(num_i[26]), .Z(n575) );
  IVSVTX2 U292 ( .A(n480), .Z(n426) );
  IVSVTX2 U293 ( .A(num_i[31]), .Z(n535) );
  ND2SVTX6 U294 ( .A(n509), .B(n508), .Z(n624) );
  CTIVSVTX2 U295 ( .A(n413), .Z(n179) );
  ND3SVTX6 U296 ( .A(n388), .B(n509), .C(n503), .Z(n299) );
  ND2SVTX4 U297 ( .A(n200), .B(n193), .Z(n537) );
  NR2SVTX4 U298 ( .A(num_i[31]), .B(num_i[27]), .Z(n238) );
  ND3ABSVTX4 U299 ( .A(num_i[12]), .B(n180), .C(n510), .Z(n412) );
  IVSVTX0H U300 ( .A(num_i[1]), .Z(n527) );
  BFSVTX2 U301 ( .A(num_i[30]), .Z(n167) );
  NR2SVTX2 U302 ( .A(num_i[20]), .B(num_i[21]), .Z(n264) );
  NR2SVTX4 U303 ( .A(num_i[15]), .B(num_i[13]), .Z(n362) );
  IVSVTX8 U304 ( .A(num_i[28]), .Z(n193) );
  IVSVTX6 U305 ( .A(num_i[30]), .Z(n200) );
  ND2SVTX6 U306 ( .A(n398), .B(n397), .Z(n410) );
  CTBUFSVTX4 U307 ( .A(num_i[19]), .Z(n589) );
  B_ND2SVTX2 U308 ( .A(n505), .B(n506), .Z(n225) );
  NR2SVTX4 U309 ( .A(num_i[20]), .B(num_i[21]), .Z(n297) );
  BFSVTX6 U310 ( .A(num_i[6]), .Z(n206) );
  IVSVTX4 U311 ( .A(num_i[5]), .Z(n180) );
  AO6ABSVTX8 U312 ( .A(n404), .B(n280), .C(n174), .Z(n401) );
  NR2SVTX8 U313 ( .A(num_i[28]), .B(num_i[30]), .Z(n365) );
  NR2SVTX8 U314 ( .A(num_i[22]), .B(num_i[23]), .Z(n510) );
  ND2SVTX8 U315 ( .A(n350), .B(n231), .Z(n358) );
  NR3ABSVTX8 U316 ( .A(n200), .B(n194), .C(n352), .Z(n530) );
  ND2ASVTX8 U317 ( .A(n232), .B(n253), .Z(n368) );
  ND3SVTX8 U318 ( .A(n210), .B(n168), .C(n332), .Z(n372) );
  ND3SVTX6 U319 ( .A(n286), .B(n642), .C(n628), .Z(n168) );
  ND2SVTX4 U320 ( .A(n169), .B(n270), .Z(n271) );
  IVSVTX4 U321 ( .A(n548), .Z(n169) );
  ND2ASVTX8 U322 ( .A(n626), .B(n276), .Z(n320) );
  AO6SVTX6 U323 ( .A(n639), .B(n325), .C(n254), .Z(n370) );
  NR2SVTX8 U324 ( .A(n249), .B(n250), .Z(n248) );
  IVSVTX12 U325 ( .A(n235), .Z(n467) );
  BFSVTX10 U326 ( .A(n636), .Z(n227) );
  IVSVTX6 U327 ( .A(n615), .Z(n197) );
  ND3SVTX6 U328 ( .A(n518), .B(n517), .C(n532), .Z(n519) );
  BFSVTX10 U329 ( .A(n601), .Z(n276) );
  ND3SVTX8 U330 ( .A(n358), .B(n170), .C(n183), .Z(n521) );
  ND3SVTX6 U331 ( .A(n448), .B(n446), .C(n507), .Z(n170) );
  AO7SVTX8 U332 ( .A(n477), .B(n460), .C(n190), .Z(n439) );
  NR2SVTX6 U333 ( .A(num_i[22]), .B(num_i[23]), .Z(n525) );
  IVSVTX6 U334 ( .A(n520), .Z(n285) );
  NR2SVTX8 U335 ( .A(n725), .B(n726), .Z(n629) );
  ND3SVTX8 U336 ( .A(n286), .B(n276), .C(n686), .Z(n700) );
  IVSVTX10 U337 ( .A(n275), .Z(n636) );
  ND3SVTX8 U338 ( .A(n697), .B(n312), .C(n368), .Z(n375) );
  AO4SVTX8 U339 ( .A(n376), .B(n375), .C(n312), .D(n695), .Z(n374) );
  ND3SVTX8 U340 ( .A(n253), .B(n171), .C(n642), .Z(n742) );
  AO1ASVTX4 U341 ( .A(num_i[4]), .B(n467), .C(n274), .D(n444), .Z(n747) );
  AO4SVTX6 U342 ( .A(n368), .B(n189), .C(n409), .D(n450), .Z(n449) );
  IVSVTX4 U343 ( .A(n319), .Z(n311) );
  ND2SVTX6 U344 ( .A(n313), .B(n372), .Z(n329) );
  ND2SVTX6 U345 ( .A(n181), .B(n687), .Z(n603) );
  ND2SVTX8 U346 ( .A(n633), .B(n634), .Z(n635) );
  AO21SVTX8 U347 ( .A(n677), .B(n678), .C(n209), .D(n227), .Z(n679) );
  ND3ABSVTX8 U348 ( .A(n428), .B(n623), .C(n732), .Z(n369) );
  MUX21NSVTX6 U349 ( .A(n639), .B(n738), .S(n363), .Z(n382) );
  AO4SVTX8 U350 ( .A(n367), .B(n216), .C(rslt_o[29]), .D(n623), .Z(n366) );
  CTBUFSVTX8 U351 ( .A(n319), .Z(n280) );
  IVSVTX12 U352 ( .A(n385), .Z(n464) );
  NR3ABSVTX8 U353 ( .A(n510), .B(n480), .C(n299), .Z(n301) );
  IVSVTX10 U354 ( .A(rslt_o[29]), .Z(n216) );
  AO6ABSVTX8 U355 ( .A(n189), .B(n283), .C(n337), .Z(n336) );
  IVSVTX8 U356 ( .A(n310), .Z(n409) );
  IVSVTX8 U357 ( .A(n640), .Z(n682) );
  ND2SVTX6 U358 ( .A(n519), .B(n539), .Z(n520) );
  IVSVTX10 U359 ( .A(n189), .Z(n313) );
  IVSVTX8 U360 ( .A(n288), .Z(n273) );
  ND2SVTX4 U361 ( .A(n650), .B(n227), .Z(n653) );
  AO7SVTX6 U362 ( .A(n546), .B(n548), .C(n198), .Z(n428) );
  IVSVTX8 U363 ( .A(n189), .Z(n188) );
  IVSVTX6 U364 ( .A(n322), .Z(n395) );
  IVSVTX8 U365 ( .A(n395), .Z(n587) );
  IVSVTX4 U366 ( .A(n402), .Z(n174) );
  ND3ABSVTX8 U367 ( .A(num_i[13]), .B(num_i[15]), .C(n433), .Z(n514) );
  IVSVTX6 U368 ( .A(n232), .Z(n608) );
  ND2SVTX4 U369 ( .A(n175), .B(n255), .Z(n256) );
  ND3SVTX6 U370 ( .A(n254), .B(n259), .C(n260), .Z(n175) );
  AO7ABSVTX4 U371 ( .A(n177), .B(n607), .C(n559), .Z(n686) );
  NR2SVTX4 U372 ( .A(n202), .B(n455), .Z(n177) );
  IVSVTX4 U373 ( .A(n288), .Z(n294) );
  ND2SVTX6 U374 ( .A(n510), .B(n388), .Z(n307) );
  NR3SVTX8 U375 ( .A(n179), .B(n178), .C(n538), .Z(n517) );
  NR2SVTX4 U376 ( .A(n206), .B(n414), .Z(n178) );
  IVSVTX4 U377 ( .A(n243), .Z(n181) );
  NR2SVTX4 U378 ( .A(n181), .B(n629), .Z(n371) );
  AO4SVTX8 U379 ( .A(n287), .B(n421), .C(n627), .D(n276), .Z(n726) );
  ND2SVTX4 U380 ( .A(n308), .B(n306), .Z(n183) );
  OR2SVTX4 U381 ( .A(num_i[24]), .B(num_i[29]), .Z(n226) );
  ND2SVTX4 U382 ( .A(n591), .B(n389), .Z(n267) );
  AO7ABSVTX6 U383 ( .A(n287), .B(n630), .C(n369), .Z(n360) );
  IVSVTX4 U384 ( .A(n621), .Z(n429) );
  IVSVTX10 U385 ( .A(num_i[29]), .Z(n194) );
  IVSVTX4 U386 ( .A(n185), .Z(n460) );
  ND2SVTX4 U387 ( .A(n716), .B(n288), .Z(n185) );
  F_ND2ASVTX2 U388 ( .A(n202), .B(n475), .Z(n712) );
  IVSVTX2 U389 ( .A(n513), .Z(n507) );
  IVSVTX2 U390 ( .A(num_i[7]), .Z(n203) );
  CTIVSVTX8 U391 ( .A(n415), .Z(keyvalues_m1[1]) );
  AN2SVTX4 U392 ( .A(n293), .B(n638), .Z(n186) );
  IVSVTX4 U393 ( .A(n341), .Z(n340) );
  AN2SVTX4 U394 ( .A(n693), .B(n391), .Z(n187) );
  ND2SVTX4 U395 ( .A(n293), .B(n379), .Z(n257) );
  IVSVTX12 U396 ( .A(n453), .Z(n470) );
  IVSVTX4 U397 ( .A(n726), .Z(n394) );
  ND3ABSVTX6 U398 ( .A(n531), .B(n307), .C(n198), .Z(n290) );
  IVSVTX8 U399 ( .A(n328), .Z(n462) );
  ND4SVTX8 U400 ( .A(n499), .B(n501), .C(n502), .D(n500), .Z(n443) );
  ND3SVTX8 U401 ( .A(n330), .B(n331), .C(n329), .Z(n328) );
  ND4SVTX8 U402 ( .A(n238), .B(n239), .C(n240), .D(n365), .Z(n364) );
  AO7SVTX4 U403 ( .A(n167), .B(n182), .C(n535), .Z(n355) );
  ND2SVTX6 U404 ( .A(n606), .B(n636), .Z(n640) );
  CTBUFSVTX4 U405 ( .A(n693), .Z(n223) );
  ND2ASVTX4 U406 ( .A(n588), .B(n425), .Z(n625) );
  AO7ABSVTX2 U407 ( .A(num_i[5]), .B(n198), .C(n592), .Z(n486) );
  F_ND2SVTX1 U408 ( .A(n673), .B(n454), .Z(n674) );
  NR2SVTX2 U409 ( .A(n705), .B(n425), .Z(n599) );
  NR2SVTX2 U410 ( .A(n622), .B(n709), .Z(n431) );
  AN2SVTX4 U411 ( .A(n591), .B(n599), .Z(n620) );
  NR2SVTX2 U412 ( .A(num_i[14]), .B(n195), .Z(n347) );
  AO3SVTX2 U413 ( .A(n676), .B(n705), .C(n675), .D(n674), .Z(n677) );
  AO7SVTX4 U414 ( .A(n720), .B(n327), .C(n719), .Z(n748) );
  IVSVTX8 U415 ( .A(n188), .Z(n191) );
  F_ND2ASVTX2 U416 ( .A(n712), .B(n484), .Z(n295) );
  IVSVTX12 U417 ( .A(n636), .Z(n189) );
  NR2SVTX6 U418 ( .A(n291), .B(n322), .Z(n275) );
  CTIVSVTX4 U419 ( .A(n278), .Z(n611) );
  CTIVSVTX2 U420 ( .A(n586), .Z(n622) );
  AO7SVTX2 U421 ( .A(num_i[2]), .B(n527), .C(n204), .Z(n529) );
  IVSVTX4 U422 ( .A(n320), .Z(n725) );
  AO1ASVTX4 U423 ( .A(n199), .B(n671), .C(n670), .D(n669), .Z(n721) );
  IVSVTX12 U424 ( .A(n467), .Z(n190) );
  IVSVTX2 U425 ( .A(n676), .Z(n671) );
  NR2SVTX2 U426 ( .A(n563), .B(n564), .Z(n656) );
  NR2SVTX6 U427 ( .A(n291), .B(n322), .Z(n235) );
  AO7SVTX4 U428 ( .A(n204), .B(n709), .C(n707), .Z(n713) );
  ND2ASVTX4 U429 ( .A(n204), .B(n454), .Z(n442) );
  IVSVTX2 U430 ( .A(n410), .Z(n547) );
  CTBUFSVTX2 U431 ( .A(num_i[14]), .Z(n673) );
  AO7SVTX4 U432 ( .A(n748), .B(n282), .C(n262), .Z(n302) );
  NR2SVTX6 U433 ( .A(n371), .B(n370), .Z(n458) );
  ND3ABSVTX4 U434 ( .A(n181), .B(n294), .C(n341), .Z(n339) );
  IVSVTX4 U435 ( .A(n741), .Z(n649) );
  IVSVTX8 U436 ( .A(n373), .Z(rslt_o[27]) );
  IVSVTX4 U437 ( .A(n326), .Z(n652) );
  AO7SVTX4 U438 ( .A(n662), .B(n409), .C(n384), .Z(n663) );
  F_ND2ASVTX2 U439 ( .A(n479), .B(n420), .Z(n646) );
  AO7SVTX6 U440 ( .A(n709), .B(n203), .C(n490), .Z(n728) );
  ND2ASVTX6 U441 ( .A(n237), .B(n583), .Z(n606) );
  IVSVTX4 U442 ( .A(n656), .Z(n648) );
  AO7NSVTX4 U443 ( .A(n202), .B(n676), .C(n661), .Z(n662) );
  ND2ASVTX4 U444 ( .A(n229), .B(n266), .Z(n583) );
  IVSVTX2 U445 ( .A(n718), .Z(n196) );
  AO7ASVTX6 U446 ( .A(n429), .B(n620), .C(n428), .Z(n430) );
  NR3ABSVTX6 U447 ( .A(num_i[4]), .B(n598), .C(n597), .Z(n610) );
  NR2ASVTX4 U448 ( .A(n673), .B(n598), .Z(n621) );
  B_ND2SVTX2 U449 ( .A(n218), .B(n454), .Z(n658) );
  ND3ASVTX2 U450 ( .A(num_i[23]), .B(n437), .C(n198), .Z(n434) );
  CTIVSVTX4 U451 ( .A(n435), .Z(n269) );
  IVSVTX8 U452 ( .A(n419), .Z(n454) );
  ND3SVTX4 U453 ( .A(n529), .B(n528), .C(n547), .Z(n400) );
  NR2SVTX2 U454 ( .A(n515), .B(n514), .Z(n518) );
  IVSVTX4 U455 ( .A(n496), .Z(n494) );
  NR3ABSVTX6 U456 ( .A(n469), .B(n535), .C(n226), .Z(n233) );
  NR2SVTX6 U457 ( .A(num_i[24]), .B(num_i[25]), .Z(n503) );
  CTBUFSVTX4 U458 ( .A(num_i[17]), .Z(n560) );
  NR2SVTX4 U459 ( .A(num_i[5]), .B(num_i[4]), .Z(n414) );
  IVSVTX6 U460 ( .A(n201), .Z(n192) );
  CTBUFSVTX2 U461 ( .A(num_i[13]), .Z(n218) );
  IVSVTX4 U462 ( .A(num_i[13]), .Z(n195) );
  AO7SVTX8 U463 ( .A(n750), .B(n262), .C(n302), .Z(keyvalues_m1[26]) );
  AO7SVTX8 U464 ( .A(rslt_o[27]), .B(n750), .C(n679), .Z(keyvalues_m1[27]) );
  NR3SVTX6 U465 ( .A(n653), .B(n652), .C(n651), .Z(n654) );
  ND2SVTX6 U466 ( .A(n406), .B(n401), .Z(n733) );
  ND3SVTX4 U467 ( .A(n310), .B(n736), .C(n440), .Z(n315) );
  AO7SVTX6 U468 ( .A(n190), .B(n461), .C(n439), .Z(keyvalues_m1[4]) );
  IVSVTX2 U469 ( .A(n478), .Z(n281) );
  IVSVTX6 U470 ( .A(n360), .Z(n325) );
  IVSVTX2 U471 ( .A(n609), .Z(n376) );
  ND2SVTX4 U472 ( .A(n648), .B(n693), .Z(n384) );
  IVSVTX2 U473 ( .A(n553), .Z(n554) );
  AO7SVTX4 U474 ( .A(n644), .B(n645), .C(n484), .Z(n420) );
  ND3SVTX4 U475 ( .A(n484), .B(n645), .C(n607), .Z(n343) );
  AO7SVTX6 U476 ( .A(n489), .B(n488), .C(n428), .Z(n490) );
  IVSVTX12 U477 ( .A(n243), .Z(n363) );
  NR2SVTX2 U478 ( .A(n660), .B(n659), .Z(n661) );
  ND2SVTX6 U479 ( .A(n266), .B(n569), .Z(n422) );
  BFSVTX2 U480 ( .A(n680), .Z(rslt_o[30]) );
  ND2ASVTX8 U481 ( .A(n593), .B(n592), .Z(n638) );
  OR2SVTX4 U482 ( .A(n334), .B(n434), .Z(n541) );
  AO7SVTX4 U483 ( .A(n668), .B(n455), .C(n335), .Z(n692) );
  IVSVTX8 U484 ( .A(n274), .Z(n222) );
  IVSVTX2 U485 ( .A(n442), .Z(n590) );
  B_ND2SVTX2 U486 ( .A(n658), .B(n182), .Z(n660) );
  ND2SVTX4 U487 ( .A(n574), .B(n269), .Z(n585) );
  NR2SVTX6 U488 ( .A(n443), .B(n521), .Z(n284) );
  IVSVTX8 U489 ( .A(n454), .Z(n455) );
  B_ND2SVTX2 U490 ( .A(num_i[8]), .B(n643), .Z(n706) );
  IVSVTX4 U491 ( .A(n437), .Z(n272) );
  NR2SVTX4 U492 ( .A(n348), .B(n346), .Z(n251) );
  ND2SVTX4 U493 ( .A(n546), .B(n436), .Z(n270) );
  B_ND2SVTX2 U494 ( .A(num_i[7]), .B(n643), .Z(n707) );
  NR2SVTX4 U495 ( .A(n476), .B(n530), .Z(n501) );
  NR3SVTX4 U496 ( .A(num_i[16]), .B(n560), .C(n351), .Z(n350) );
  NR2SVTX6 U497 ( .A(num_i[16]), .B(num_i[17]), .Z(n509) );
  CTIVSVTX2 U498 ( .A(num_i[4]), .Z(n199) );
  NR2SVTX4 U499 ( .A(num_i[9]), .B(num_i[8]), .Z(n397) );
  CTBUFSVTX12 U500 ( .A(num_i[11]), .Z(n552) );
  NR2SVTX4 U501 ( .A(num_i[9]), .B(num_i[8]), .Z(n413) );
  NR2SVTX6 U502 ( .A(num_i[29]), .B(num_i[25]), .Z(n289) );
  IVSVTX4 U503 ( .A(num_i[21]), .Z(n201) );
  CTIVSVTX4 U504 ( .A(num_i[3]), .Z(n204) );
  ND3ABSVTX8 U505 ( .A(n205), .B(n187), .C(n374), .Z(keyvalues_m1[20]) );
  NR2SVTX4 U506 ( .A(n327), .B(n640), .Z(n205) );
  CTBUFSVTX8 U507 ( .A(n683), .Z(n219) );
  AO2SVTX8 U508 ( .A(n692), .B(n691), .C(n717), .D(n683), .Z(n283) );
  AO7ABSVTX8 U509 ( .A(n613), .B(n628), .C(n317), .Z(n737) );
  ND2SVTX4 U510 ( .A(n259), .B(n260), .Z(n687) );
  AO2SVTX8 U511 ( .A(n280), .B(n261), .C(n311), .D(n608), .Z(n260) );
  IVSVTX6 U512 ( .A(n190), .Z(n215) );
  ND3SVTX8 U513 ( .A(n451), .B(n191), .C(n283), .Z(n217) );
  NR2SVTX6 U514 ( .A(num_i[28]), .B(num_i[30]), .Z(n452) );
  ND2SVTX6 U515 ( .A(n642), .B(n258), .Z(n699) );
  ND2SVTX8 U516 ( .A(n297), .B(n525), .Z(n538) );
  ND2SVTX6 U517 ( .A(n377), .B(n378), .Z(n739) );
  IVSVTX4 U518 ( .A(n456), .Z(n207) );
  AO2SVTX6 U519 ( .A(n494), .B(n493), .C(n207), .D(n575), .Z(n500) );
  IVSVTX12 U520 ( .A(n319), .Z(n288) );
  NR2SVTX4 U521 ( .A(n628), .B(n721), .Z(n209) );
  ND2SVTX4 U522 ( .A(n196), .B(n691), .Z(n579) );
  OR2ABSVTX8 U523 ( .A(num_i[23]), .B(n389), .Z(n244) );
  ND3ASVTX6 U524 ( .A(num_i[27]), .B(n562), .C(n193), .Z(n234) );
  ND2ASVTX8 U525 ( .A(n189), .B(n737), .Z(n316) );
  IVSVTX4 U526 ( .A(n212), .Z(n310) );
  ND2SVTX2 U527 ( .A(n224), .B(n601), .Z(n212) );
  ND2SVTX4 U528 ( .A(n213), .B(n214), .Z(n453) );
  ND2SVTX4 U529 ( .A(n190), .B(n734), .Z(n213) );
  ND2SVTX4 U530 ( .A(n309), .B(n215), .Z(n214) );
  NR3ABSVTX2 U531 ( .A(n475), .B(num_i[4]), .C(n216), .Z(n478) );
  ND3SVTX8 U532 ( .A(n316), .B(n315), .C(n314), .Z(keyvalues_m1[15]) );
  BFSVTX2 U533 ( .A(num_i[15]), .Z(n230) );
  NR2ASVTX6 U534 ( .A(n181), .B(n748), .Z(n724) );
  ND2SVTX2 U535 ( .A(n323), .B(n224), .Z(n740) );
  AN2SVTX4 U536 ( .A(n464), .B(n601), .Z(n693) );
  AO7SVTX6 U537 ( .A(n743), .B(n744), .C(n217), .Z(n745) );
  IVSVTX12 U538 ( .A(n287), .Z(n732) );
  ND2ASVTX8 U539 ( .A(num_i[25]), .B(n511), .Z(n531) );
  IVSVTX8 U540 ( .A(num_i[25]), .Z(n562) );
  BFSVTX4 U541 ( .A(n548), .Z(n435) );
  ND3SVTX6 U542 ( .A(n637), .B(n416), .C(n319), .Z(n377) );
  NR3ASVTX6 U543 ( .A(rslt_o[29]), .B(n551), .C(n550), .Z(n557) );
  NR2SVTX4 U544 ( .A(n410), .B(n528), .Z(n481) );
  NR4SVTX8 U545 ( .A(num_i[7]), .B(num_i[6]), .C(num_i[5]), .D(num_i[4]), .Z(
        n528) );
  ND2SVTX4 U546 ( .A(n262), .B(n701), .Z(n702) );
  AO7SVTX8 U547 ( .A(n442), .B(n197), .C(n441), .Z(n642) );
  IVSVTX6 U548 ( .A(n614), .Z(n367) );
  AO4SVTX8 U549 ( .A(n731), .B(n313), .C(n312), .D(n730), .Z(keyvalues_m1[8])
         );
  ND3SVTX8 U550 ( .A(n342), .B(n343), .C(n344), .Z(n341) );
  ND2SVTX6 U551 ( .A(n525), .B(n388), .Z(n361) );
  ND3ASVTX8 U552 ( .A(n570), .B(n423), .C(n422), .Z(n694) );
  BFSVTX1 U553 ( .A(n628), .Z(rslt_o[28]) );
  ND2SVTX4 U554 ( .A(n407), .B(n215), .Z(n406) );
  IVSVTX6 U555 ( .A(n363), .Z(n254) );
  ND3SVTX8 U556 ( .A(n424), .B(n604), .C(n603), .Z(keyvalues_m1[17]) );
  ND2ASVTX8 U557 ( .A(n704), .B(n379), .Z(n421) );
  IVSVTX4 U558 ( .A(n739), .Z(n221) );
  ND3ASVTX6 U559 ( .A(n622), .B(n222), .C(n428), .Z(n524) );
  ND2SVTX4 U560 ( .A(n188), .B(n359), .Z(n634) );
  AO7SVTX8 U561 ( .A(n617), .B(n657), .C(n616), .Z(n614) );
  NR2SVTX4 U562 ( .A(n725), .B(n254), .Z(n393) );
  ND2SVTX4 U563 ( .A(n473), .B(n481), .Z(n436) );
  IVSVTX4 U564 ( .A(n225), .Z(n473) );
  AO8DSVTX6 U565 ( .A(n403), .B(n540), .C(n287), .D(n643), .Z(n402) );
  ND3ABSVTX8 U566 ( .A(n471), .B(n483), .C(n301), .Z(n437) );
  MUX21NSVTX4 U567 ( .A(n296), .B(n295), .S(n628), .Z(n457) );
  ND2SVTX4 U568 ( .A(n694), .B(n228), .Z(n259) );
  NR2ASVTX6 U569 ( .A(rslt_o[29]), .B(n287), .Z(n228) );
  AO7SVTX6 U570 ( .A(n304), .B(n400), .C(n396), .Z(n241) );
  IVSVTX4 U571 ( .A(n298), .Z(n574) );
  ND2ASVTX8 U572 ( .A(n298), .B(n561), .Z(n607) );
  NR2ASVTX6 U573 ( .A(n410), .B(n211), .Z(n549) );
  AO7ABSVTX6 U574 ( .A(n693), .B(n717), .C(n579), .Z(n651) );
  NR3ABSVTX8 U575 ( .A(n264), .B(n503), .C(n263), .Z(n231) );
  BFSVTX2 U576 ( .A(num_i[18]), .Z(n584) );
  AO17SVTX6 U577 ( .A(n552), .B(n533), .C(n399), .D(n532), .Z(n396) );
  IVSVTX2 U578 ( .A(n595), .Z(n381) );
  ND2ASVTX8 U579 ( .A(n224), .B(n614), .Z(n232) );
  NR3ABSVTX2 U580 ( .A(n475), .B(num_i[3]), .C(n287), .Z(n323) );
  AO7ASVTX6 U581 ( .A(n206), .B(n709), .C(n524), .Z(n710) );
  OR2SVTX8 U582 ( .A(n624), .B(n538), .Z(n591) );
  ND4ABSVTX4 U583 ( .A(n229), .B(n586), .C(n533), .D(n532), .Z(n534) );
  IVSVTX4 U584 ( .A(n534), .Z(n246) );
  MUX21NSVTX6 U585 ( .A(n710), .B(n711), .S(n287), .Z(n731) );
  ND2ASVTX8 U586 ( .A(n234), .B(n233), .Z(n502) );
  ND2SVTX8 U587 ( .A(n244), .B(n236), .Z(n322) );
  NR2SVTX8 U588 ( .A(n242), .B(n241), .Z(n236) );
  MUX21NSVTX8 U589 ( .A(n735), .B(n605), .S(n467), .Z(n349) );
  ND3ASVTX8 U590 ( .A(n251), .B(n245), .C(n248), .Z(n291) );
  IVSVTX4 U591 ( .A(n606), .Z(n735) );
  NR2SVTX4 U592 ( .A(n582), .B(n274), .Z(n237) );
  NR2SVTX6 U593 ( .A(num_i[24]), .B(num_i[29]), .Z(n239) );
  NR2SVTX6 U594 ( .A(num_i[26]), .B(num_i[25]), .Z(n240) );
  ND3ASVTX6 U595 ( .A(n530), .B(n303), .C(n358), .Z(n242) );
  NR2SVTX8 U596 ( .A(n322), .B(n291), .Z(n243) );
  NR2SVTX6 U597 ( .A(n247), .B(n246), .Z(n245) );
  NR2ASVTX6 U598 ( .A(n589), .B(n290), .Z(n249) );
  AO7ABSVTX8 U599 ( .A(n345), .B(n389), .C(n539), .Z(n250) );
  NR2SVTX6 U600 ( .A(n492), .B(n456), .Z(n493) );
  ND2SVTX8 U601 ( .A(n194), .B(n193), .Z(n456) );
  ND4SVTX4 U602 ( .A(n181), .B(n700), .C(n685), .D(n699), .Z(n255) );
  ND2ASVTX8 U603 ( .A(n257), .B(n273), .Z(n685) );
  ND2SVTX6 U604 ( .A(n688), .B(n256), .Z(keyvalues_m1[18]) );
  AO4SVTX6 U605 ( .A(n189), .B(n451), .C(n181), .D(n338), .Z(n337) );
  ND4SVTX6 U606 ( .A(num_i[15]), .B(n193), .C(n194), .D(n508), .Z(n263) );
  NR2SVTX8 U607 ( .A(num_i[18]), .B(num_i[19]), .Z(n508) );
  NR2SVTX8 U608 ( .A(n605), .B(n363), .Z(n391) );
  AO2SVTX8 U609 ( .A(n585), .B(n584), .C(n472), .D(n586), .Z(n605) );
  ND2SVTX4 U610 ( .A(n310), .B(n747), .Z(n415) );
  NR2SVTX6 U611 ( .A(num_i[19]), .B(num_i[16]), .Z(n505) );
  ND3ABSVTX8 U612 ( .A(n643), .B(n272), .C(n271), .Z(n385) );
  IVSVTX12 U613 ( .A(n601), .Z(n287) );
  ND2SVTX8 U614 ( .A(n285), .B(n284), .Z(n601) );
  AO7ABSVTX8 U615 ( .A(n746), .B(n391), .C(n745), .Z(keyvalues_m1[22]) );
  ND3SVTX8 U616 ( .A(n459), .B(n702), .C(n703), .Z(keyvalues_m1[19]) );
  ND2SVTX8 U617 ( .A(n690), .B(n292), .Z(keyvalues_m1[2]) );
  IVSVTX12 U618 ( .A(n601), .Z(n319) );
  ND2SVTX4 U619 ( .A(n569), .B(n475), .Z(n278) );
  IVSVTX4 U620 ( .A(n279), .Z(n335) );
  MUX21NSVTX8 U621 ( .A(n727), .B(n713), .S(n319), .Z(n309) );
  ND2SVTX4 U622 ( .A(n646), .B(n280), .Z(n741) );
  IVSVTX4 U623 ( .A(n723), .Z(n282) );
  ND2ASVTX8 U624 ( .A(n280), .B(n749), .Z(n723) );
  IVSVTX4 U625 ( .A(n416), .Z(n286) );
  MUX21NSVTX8 U626 ( .A(n711), .B(n716), .S(n287), .Z(n734) );
  NR2SVTX8 U627 ( .A(num_i[26]), .B(num_i[24]), .Z(n511) );
  ND2SVTX8 U628 ( .A(n289), .B(n511), .Z(n513) );
  ND2SVTX4 U629 ( .A(n188), .B(n457), .Z(n292) );
  AO21SVTX8 U630 ( .A(n580), .B(n652), .C(n651), .D(n312), .Z(n581) );
  NR2SVTX4 U631 ( .A(n355), .B(n354), .Z(n303) );
  ND2SVTX4 U632 ( .A(n533), .B(n532), .Z(n304) );
  ND2SVTX8 U633 ( .A(n365), .B(n305), .Z(n485) );
  NR2SVTX6 U634 ( .A(num_i[29]), .B(num_i[31]), .Z(n305) );
  AO1ABSVTX6 U635 ( .A(num_i[19]), .B(num_i[14]), .C(n307), .D(n485), .Z(n306)
         );
  AO6SVTX6 U636 ( .A(n543), .B(n624), .C(n531), .Z(n308) );
  MUX21NSVTX8 U637 ( .A(n731), .B(n309), .S(n190), .Z(n468) );
  ND2SVTX4 U638 ( .A(n366), .B(n294), .Z(n317) );
  IVSVTX12 U639 ( .A(n318), .Z(n683) );
  ND2ASVTX8 U640 ( .A(n601), .B(n484), .Z(n318) );
  MUX21NSVTX8 U641 ( .A(n710), .B(n631), .S(n288), .Z(n729) );
  AO2SVTX8 U642 ( .A(n393), .B(n394), .C(n359), .D(n312), .Z(keyvalues_m1[12])
         );
  ND2SVTX6 U643 ( .A(num_i[27]), .B(n193), .Z(n352) );
  NR3SVTX8 U644 ( .A(n382), .B(n324), .C(n380), .Z(n641) );
  NR2SVTX4 U645 ( .A(n188), .B(n325), .Z(n324) );
  ND2ASVTX8 U646 ( .A(rslt_o[29]), .B(n273), .Z(n327) );
  ND3ASVTX6 U647 ( .A(rslt_o[29]), .B(n694), .C(n273), .Z(n326) );
  IVSVTX4 U648 ( .A(n327), .Z(n746) );
  ND2SVTX4 U649 ( .A(n186), .B(n253), .Z(n332) );
  ND2ASVTX8 U650 ( .A(n381), .B(n596), .Z(n379) );
  ND2SVTX6 U651 ( .A(n686), .B(n683), .Z(n338) );
  AO7SVTX6 U652 ( .A(n273), .B(n340), .C(n338), .Z(n695) );
  ND3SVTX8 U653 ( .A(n696), .B(n339), .C(n336), .Z(keyvalues_m1[21]) );
  ND2SVTX4 U654 ( .A(n216), .B(n642), .Z(n342) );
  ND2SVTX4 U655 ( .A(n347), .B(n545), .Z(n346) );
  IVSVTX4 U656 ( .A(n544), .Z(n348) );
  ND2SVTX4 U657 ( .A(n219), .B(n349), .Z(n424) );
  ND2SVTX4 U658 ( .A(n746), .B(n349), .Z(n696) );
  AO2SVTX6 U659 ( .A(n313), .B(n698), .C(n349), .D(n223), .Z(n703) );
  ND2SVTX4 U660 ( .A(n357), .B(n200), .Z(n351) );
  NR2SVTX8 U661 ( .A(num_i[22]), .B(num_i[26]), .Z(n357) );
  MUX21NSVTX8 U662 ( .A(n631), .B(n630), .S(n732), .Z(n359) );
  NR2SVTX8 U663 ( .A(n513), .B(n386), .Z(n532) );
  ND3SVTX8 U664 ( .A(n506), .B(n505), .C(n452), .Z(n386) );
  ND4ABSVTX8 U665 ( .A(n410), .B(n203), .C(n533), .D(n532), .Z(n539) );
  NR3ABSVTX8 U666 ( .A(n362), .B(n433), .C(n361), .Z(n533) );
  NR2SVTX4 U667 ( .A(num_i[27]), .B(num_i[26]), .Z(n387) );
  ND2SVTX6 U668 ( .A(n618), .B(n619), .Z(n639) );
  ND2SVTX4 U669 ( .A(n191), .B(n372), .Z(n604) );
  ND3ABSVTX8 U670 ( .A(n484), .B(n383), .C(n311), .Z(n738) );
  NR2ASVTX6 U671 ( .A(n665), .B(n274), .Z(n570) );
  AO6SVTX2 U672 ( .A(n274), .B(n665), .C(num_i[28]), .Z(n666) );
  IVSVTX4 U673 ( .A(n386), .Z(n448) );
  IVSVTX12 U674 ( .A(n464), .Z(rslt_o[29]) );
  NR2SVTX8 U675 ( .A(num_i[21]), .B(num_i[20]), .Z(n388) );
  ND2SVTX6 U676 ( .A(n387), .B(n392), .Z(n466) );
  ND2SVTX4 U677 ( .A(n218), .B(n475), .Z(n592) );
  AO2SVTX4 U678 ( .A(n391), .B(n219), .C(n682), .D(n223), .Z(n688) );
  NR2SVTX6 U679 ( .A(num_i[25]), .B(num_i[24]), .Z(n392) );
  NR3SVTX8 U680 ( .A(n537), .B(n536), .C(n466), .Z(n545) );
  NR2SVTX6 U681 ( .A(num_i[11]), .B(num_i[10]), .Z(n398) );
  MUX21NSVTX4 U682 ( .A(n206), .B(num_i[4]), .S(n319), .Z(n407) );
  NR2ASVTX6 U683 ( .A(n204), .B(n587), .Z(n403) );
  ND3ABSVTX8 U684 ( .A(n405), .B(n587), .C(n540), .Z(n404) );
  MUX21NSVTX8 U685 ( .A(n730), .B(n729), .S(n227), .Z(keyvalues_m1[9]) );
  MUX21NSVTX8 U686 ( .A(n729), .B(n632), .S(n313), .Z(keyvalues_m1[10]) );
  IVSVTX4 U687 ( .A(num_i[24]), .Z(n482) );
  ND3SVTX6 U688 ( .A(n705), .B(n526), .C(n388), .Z(n411) );
  IVSVTX4 U689 ( .A(num_i[6]), .Z(n705) );
  IVSVTX4 U690 ( .A(n484), .Z(n416) );
  NR2ASVTX6 U691 ( .A(n429), .B(n620), .Z(n612) );
  ND2SVTX4 U692 ( .A(n545), .B(n544), .Z(n419) );
  NR2SVTX4 U693 ( .A(n624), .B(n538), .Z(n544) );
  NR2SVTX4 U694 ( .A(num_i[27]), .B(num_i[26]), .Z(n480) );
  NR2SVTX8 U695 ( .A(n277), .B(n319), .Z(n619) );
  NR2SVTX6 U696 ( .A(num_i[17]), .B(num_i[18]), .Z(n506) );
  AO6SVTX8 U697 ( .A(n549), .B(n473), .C(n548), .Z(n561) );
  IVSVTX4 U698 ( .A(n425), .Z(n598) );
  ND2SVTX4 U699 ( .A(n427), .B(n475), .Z(n708) );
  AO20SVTX8 U700 ( .A(n546), .B(n435), .C(n198), .D(n229), .Z(n427) );
  OR2SVTX8 U701 ( .A(n426), .B(n496), .Z(n548) );
  NR2SVTX4 U702 ( .A(n611), .B(n610), .Z(n623) );
  NR2SVTX4 U703 ( .A(num_i[15]), .B(num_i[14]), .Z(n526) );
  NR2SVTX6 U704 ( .A(num_i[12]), .B(num_i[14]), .Z(n433) );
  IVSVTX4 U705 ( .A(n538), .Z(n546) );
  IVSVTX4 U706 ( .A(num_i[22]), .Z(n504) );
  ND2SVTX4 U707 ( .A(n735), .B(n190), .Z(n440) );
  MUX21SVTX4 U708 ( .A(n734), .B(n461), .S(n190), .Z(n438) );
  AO2SVTX6 U709 ( .A(n472), .B(n552), .C(n475), .D(n589), .Z(n441) );
  NR2SVTX4 U710 ( .A(num_i[3]), .B(n467), .Z(n444) );
  NR4SVTX8 U711 ( .A(num_i[12]), .B(n192), .C(n665), .D(n447), .Z(n446) );
  AO7SVTX6 U712 ( .A(num_i[10]), .B(n552), .C(n195), .Z(n447) );
  IVSVTX4 U713 ( .A(n449), .Z(n459) );
  ND2SVTX4 U714 ( .A(n717), .B(n467), .Z(n450) );
  ND2SVTX4 U715 ( .A(n694), .B(n693), .Z(n451) );
  NR2SVTX2 U716 ( .A(n582), .B(n680), .Z(n564) );
  ND2SVTX4 U717 ( .A(n574), .B(n561), .Z(n680) );
  AO7SVTX6 U718 ( .A(n558), .B(n557), .C(n556), .Z(n664) );
  NR2ASVTX2 U719 ( .A(n203), .B(n484), .Z(n553) );
  ND3ABSVTX6 U720 ( .A(n498), .B(n456), .C(n497), .Z(n499) );
  ND3SVTX4 U721 ( .A(n700), .B(n685), .C(n699), .Z(n701) );
  MUX21NSVTX8 U722 ( .A(n713), .B(n714), .S(n287), .Z(n461) );
  NR2ASVTX2 U723 ( .A(num_i[7]), .B(n455), .Z(n645) );
  AO2SVTX2 U724 ( .A(n475), .B(n571), .C(n472), .D(n673), .Z(n573) );
  IVSVTX12 U725 ( .A(n462), .Z(keyvalues_m1[16]) );
  AN2SVTX4 U726 ( .A(n319), .B(n715), .Z(n477) );
  ND2ASVTX1 U727 ( .A(n594), .B(n475), .Z(n595) );
  AO7SVTX8 U728 ( .A(n373), .B(n722), .C(n581), .Z(keyvalues_m1[24]) );
  AO7ABSVTX4 U729 ( .A(n648), .B(n691), .C(n647), .Z(n743) );
  ND2SVTX2 U730 ( .A(n691), .B(n717), .Z(n609) );
  IVSVTX2 U731 ( .A(n692), .Z(n568) );
  IVSVTX2 U732 ( .A(num_i[20]), .Z(n495) );
  NR3SVTX2 U733 ( .A(num_i[6]), .B(num_i[2]), .C(num_i[3]), .Z(n515) );
  AN2ABSVTX8 U734 ( .A(n312), .B(n740), .Z(keyvalues_m1[0]) );
  IVSVTX12 U735 ( .A(n458), .Z(n465) );
  AO6ASVTX8 U736 ( .A(n253), .B(n664), .C(n567), .Z(n722) );
  ND2SVTX4 U737 ( .A(n189), .B(n632), .Z(n633) );
  MUX21NSVTX6 U738 ( .A(n728), .B(n727), .S(n319), .Z(n730) );
  ND3ASVTX4 U739 ( .A(n705), .B(n680), .C(n454), .Z(n572) );
  IVSVTX4 U740 ( .A(n504), .Z(n469) );
  IVSVTX4 U741 ( .A(n697), .Z(n698) );
  IVSVTX4 U742 ( .A(n597), .Z(n600) );
  NR2SVTX2 U743 ( .A(rslt_o[29]), .B(n718), .Z(n678) );
  AO7SVTX6 U744 ( .A(n709), .B(n668), .C(n523), .Z(n631) );
  ND2SVTX4 U745 ( .A(n694), .B(n683), .Z(n697) );
  NR2ASVTX2 U746 ( .A(n192), .B(n680), .Z(n659) );
  ND2SVTX4 U747 ( .A(n683), .B(n196), .Z(n719) );
  NR2ASVTX6 U748 ( .A(n201), .B(n496), .Z(n497) );
  ND2ASVTX8 U749 ( .A(n487), .B(n198), .Z(n709) );
  IVSVTX10 U750 ( .A(n641), .Z(keyvalues_m1[14]) );
  NR2SVTX2 U751 ( .A(n612), .B(n484), .Z(n613) );
  AO6CSVTX2 U752 ( .A(n484), .B(n588), .C(n454), .Z(n555) );
  AO2ABSVTX4 U753 ( .C(n428), .D(n486), .A(n709), .B(n229), .Z(n627) );
  AO2SVTX4 U754 ( .A(n222), .B(n192), .C(n472), .D(n218), .Z(n559) );
  ND2SVTX2 U755 ( .A(n605), .B(n467), .Z(n736) );
  AN2SVTX0H U756 ( .A(num_i[3]), .B(n624), .Z(n474) );
  IVSVTX2 U757 ( .A(num_i[23]), .Z(n492) );
  AN2SVTX0H U758 ( .A(num_i[23]), .B(n643), .Z(n479) );
  AO7SVTX2 U759 ( .A(n617), .B(n197), .C(n616), .Z(n618) );
  ND2SVTX8 U760 ( .A(n562), .B(n482), .Z(n496) );
  IVSVTX4 U761 ( .A(n625), .Z(n489) );
  BFSVTX6 U762 ( .A(num_i[20]), .Z(n665) );
  IVSVTX4 U763 ( .A(n589), .Z(n543) );
  ND2SVTX4 U764 ( .A(n535), .B(n194), .Z(n536) );
  NR2SVTX4 U765 ( .A(n644), .B(n541), .Z(n558) );
  IVSVTX0H U766 ( .A(num_i[27]), .Z(n542) );
  ND2SVTX4 U767 ( .A(n574), .B(n561), .Z(n615) );
  NR2ASVTX2 U768 ( .A(n590), .B(n615), .Z(n550) );
  ND2SVTX4 U769 ( .A(n555), .B(n554), .Z(n556) );
  AO7SVTX2 U770 ( .A(n229), .B(n455), .C(n562), .Z(n563) );
  IVSVTX4 U771 ( .A(n650), .Z(n580) );
  IVSVTX0H U772 ( .A(n575), .Z(n576) );
  AO7SVTX2 U773 ( .A(n622), .B(n455), .C(n576), .Z(n577) );
  AO6ABSVTX4 U774 ( .A(n578), .B(n585), .C(n577), .Z(n718) );
  NR2SVTX8 U775 ( .A(n293), .B(n287), .Z(n691) );
  AO7ABSVTX4 U776 ( .A(n598), .B(n474), .C(n625), .Z(n637) );
  NR2SVTX8 U777 ( .A(n654), .B(n655), .Z(keyvalues_m1[23]) );
  AO20SVTX4 U778 ( .A(n668), .B(rslt_o[29]), .C(n667), .D(n455), .Z(n669) );
  NR2SVTX2 U779 ( .A(n167), .B(n672), .Z(n675) );
  NR2ASVTX1 U780 ( .A(num_i[3]), .B(n198), .Z(n689) );
  NR3SVTX8 U781 ( .A(n705), .B(n274), .C(n704), .Z(n716) );
  AO7SVTX4 U782 ( .A(n709), .B(n202), .C(n708), .Z(n727) );
  NR2ASVTX2 U783 ( .A(n643), .B(n712), .Z(n714) );
  NR2ASVTX1 U784 ( .A(num_i[4]), .B(n198), .Z(n715) );
  IVSVTX2 U785 ( .A(n717), .Z(n720) );
  IVSVTX4 U786 ( .A(n721), .Z(n749) );
  AO2ASVTX8 U787 ( .C(n724), .D(n723), .A(rslt_o[27]), .B(n722), .Z(
        keyvalues_m1[25]) );
  IVSVTX12 U788 ( .A(n733), .Z(keyvalues_m1[3]) );
endmodule

