
module m_rangemapping ( N, O );
  input [31:0] N;
  output [31:0] O;
  wire   n211, n212, n213, n214, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n263, n264, n265, n266, n267, n268,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n324, n325, n326,
         n327, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n505, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n719, n720, n721, n722, n723, n724,
         n725, n726, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n915, n917, n918, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814;

  F_ENSVTX2 U296 ( .A(n245), .B(n1748), .Z(O[17]) );
  IVSVTX0H U297 ( .A(n1329), .Z(O[30]) );
  EOSVTX1 U298 ( .A(n1763), .B(n1762), .Z(O[10]) );
  EOSVTX1 U299 ( .A(n1786), .B(n1785), .Z(O[7]) );
  EOSVTX0H U300 ( .A(n1777), .B(n1776), .Z(O[3]) );
  EOSVTX0H U301 ( .A(n1767), .B(n1766), .Z(O[9]) );
  ENSVTX0H U302 ( .A(n1771), .B(n1770), .Z(O[8]) );
  IVSVTX12 U303 ( .A(n1285), .Z(O[31]) );
  ENSVTX1 U304 ( .A(n1696), .B(n1695), .Z(O[13]) );
  ENSVTX1 U305 ( .A(n1272), .B(n1271), .Z(O[11]) );
  ENSVTX0H U306 ( .A(n1789), .B(n1788), .Z(O[1]) );
  ENSVTX1 U307 ( .A(n1700), .B(n1753), .Z(O[12]) );
  ENSVTX0H U308 ( .A(n1715), .B(n1784), .Z(O[6]) );
  ENSVTX0H U309 ( .A(n1795), .B(n1794), .Z(O[5]) );
  BFSVTX2 U310 ( .A(n1642), .Z(n403) );
  AO6SVTX1 U311 ( .A(n1770), .B(n1769), .C(n230), .Z(n1766) );
  AO6SVTX1 U312 ( .A(n1788), .B(n1787), .C(n1708), .Z(n1709) );
  AO7SVTX1 U313 ( .A(n1762), .B(n1270), .C(n1438), .Z(n1271) );
  IVSVTX0H U314 ( .A(n1699), .Z(n1753) );
  AO7SVTX1 U315 ( .A(n1793), .B(n1798), .C(n1796), .Z(n1794) );
  AO7SVTX1 U316 ( .A(n1694), .B(n1699), .C(n1697), .Z(n1695) );
  F_ND2SVTX0H U317 ( .A(n1703), .B(n1702), .Z(n1710) );
  F_ND2SVTX0H U318 ( .A(n694), .B(n1778), .Z(n1779) );
  IVSVTX0H U319 ( .A(n1725), .Z(n1682) );
  IVSVTX0H U320 ( .A(n1701), .Z(n1702) );
  IVSVTX0H U321 ( .A(n702), .Z(n1438) );
  AO6SVTX1 U322 ( .A(n1770), .B(n1266), .C(n721), .Z(n1762) );
  IVSVTX0H U323 ( .A(n1802), .Z(n1804) );
  BFSVTX2 U324 ( .A(n461), .Z(n320) );
  IVSVTX2 U325 ( .A(n707), .Z(n708) );
  F_ND2SVTX1 U326 ( .A(n429), .B(n430), .Z(n1747) );
  CTIVSVTX2 U327 ( .A(n1684), .Z(n223) );
  IVSVTX0H U328 ( .A(n1761), .Z(n1270) );
  IVSVTX0H U329 ( .A(n1797), .Z(n1793) );
  IVSVTX0H U330 ( .A(n1755), .Z(n1756) );
  IVSVTX0H U331 ( .A(n1783), .Z(n751) );
  IVSVTX0H U332 ( .A(n347), .Z(n1708) );
  NR2SVTX2 U333 ( .A(n1722), .B(n1683), .Z(n1686) );
  IVSVTX0H U334 ( .A(n1698), .Z(n1694) );
  AN2SVTX2 U335 ( .A(n1809), .B(n352), .Z(n794) );
  AO7SVTX1 U336 ( .A(n1714), .B(n1798), .C(n1713), .Z(n1784) );
  BFSVTX0H U337 ( .A(n1792), .Z(n1796) );
  IVSVTX6 U338 ( .A(n487), .Z(n782) );
  CTIVSVTX2 U339 ( .A(n1739), .Z(n707) );
  IVSVTX0H U340 ( .A(n1782), .Z(n1783) );
  IVSVTX0H U341 ( .A(n1434), .Z(n1266) );
  IVSVTX0H U342 ( .A(n1712), .Z(n1713) );
  BFSVTX0H U343 ( .A(n1704), .Z(n1802) );
  AO7SVTX1 U344 ( .A(n753), .B(n765), .C(n1808), .Z(n1810) );
  AO6NSVTX1 U345 ( .A(n230), .B(n238), .C(n1265), .Z(n721) );
  ND3SVTX2 U346 ( .A(n409), .B(n354), .C(n353), .Z(n1809) );
  BFSVTX0H U347 ( .A(n349), .Z(n347) );
  BFSVTX0H U348 ( .A(n1437), .Z(n1761) );
  ND2ASVTX1 U349 ( .A(n1496), .B(n1754), .Z(n1755) );
  BFSVTX0H U350 ( .A(n756), .Z(n238) );
  BFSVTX0H U351 ( .A(n1765), .Z(n230) );
  IVSVTX6 U352 ( .A(n1683), .Z(n286) );
  IVSVTX4 U353 ( .A(n1735), .Z(n731) );
  BFSVTX2 U354 ( .A(n383), .Z(n409) );
  ND2ASVTX6 U355 ( .A(n1667), .B(n1666), .Z(n1670) );
  IVSVTX0H U356 ( .A(n1436), .Z(n367) );
  NR2SVTX6 U357 ( .A(n1641), .B(n544), .Z(n1735) );
  ND2SVTX6 U358 ( .A(n1639), .B(n1640), .Z(n438) );
  NR2SVTX6 U359 ( .A(n1681), .B(n1680), .Z(n1725) );
  AO7ABSVTX2 U360 ( .A(n279), .B(n456), .C(n213), .Z(n455) );
  IVSVTX6 U361 ( .A(n1716), .Z(n765) );
  IVSVTX4 U362 ( .A(n445), .Z(n394) );
  IVSVTX0H U363 ( .A(n1719), .Z(n456) );
  CTIVSVTX4 U364 ( .A(n1669), .Z(n1663) );
  IVSVTX0H U365 ( .A(n1637), .Z(n281) );
  IVSVTX4 U366 ( .A(n1664), .Z(n1657) );
  ND3SVTX6 U367 ( .A(n771), .B(n380), .C(n379), .Z(n1746) );
  AO6SVTX4 U368 ( .A(n443), .B(n523), .C(n771), .Z(n430) );
  ND2ASVTX4 U369 ( .A(n1161), .B(n287), .Z(n429) );
  IVSVTX0H U370 ( .A(n1674), .Z(n1600) );
  F_ENSVTX2 U371 ( .A(n1581), .B(n1583), .Z(n771) );
  NR2SVTX2 U372 ( .A(n431), .B(n443), .Z(n1745) );
  IVSVTX2 U373 ( .A(n1582), .Z(n523) );
  AO7ASVTX6 U374 ( .A(n534), .B(n545), .C(n532), .Z(n1667) );
  ND3SVTX4 U375 ( .A(n383), .B(n293), .C(n764), .Z(n258) );
  ENSVTX1 U376 ( .A(n1659), .B(n1658), .Z(n1653) );
  IVSVTX0H U377 ( .A(n1636), .Z(n433) );
  IVSVTX0H U378 ( .A(n1591), .Z(n1592) );
  AO7SVTX6 U379 ( .A(n543), .B(n1716), .C(n1617), .Z(n391) );
  AO6NSVTX1 U380 ( .A(n1570), .B(n464), .C(n1564), .Z(n711) );
  ND2ASVTX4 U381 ( .A(n510), .B(n383), .Z(n1582) );
  ENSVTX0H U382 ( .A(n1585), .B(n1586), .Z(n1581) );
  IVSVTX6 U383 ( .A(n443), .Z(n287) );
  BFSVTX6 U384 ( .A(n1656), .Z(n224) );
  IVSVTX0H U385 ( .A(n1617), .Z(n510) );
  BFSVTX1 U386 ( .A(n1676), .Z(n755) );
  F_ND2ASVTX2 U387 ( .A(n1402), .B(n1718), .Z(n221) );
  IVSVTX2 U388 ( .A(n543), .Z(n240) );
  IVSVTX0H U389 ( .A(n1632), .Z(n220) );
  IVSVTX0H U390 ( .A(n1563), .Z(n1386) );
  HA1SVTX2 U391 ( .A(n1650), .B(n738), .CO(n1602), .S(n1659) );
  BFSVTX2 U392 ( .A(n1599), .Z(n1601) );
  ND3SVTX4 U393 ( .A(n1718), .B(n1631), .C(n764), .Z(n1634) );
  ND2SVTX2 U394 ( .A(n291), .B(n1574), .Z(n1679) );
  IVSVTX0H U395 ( .A(n1610), .Z(n1611) );
  IVSVTX0H U396 ( .A(n1586), .Z(n1584) );
  IVSVTX0H U397 ( .A(n1569), .Z(n1432) );
  CTBUFSVTX4 U398 ( .A(n1607), .Z(n616) );
  BFSVTX2 U399 ( .A(n1565), .Z(n464) );
  BFSVTX2 U400 ( .A(n1579), .Z(n1586) );
  IVSVTX8 U401 ( .A(n1646), .Z(n1604) );
  ND2ASVTX4 U402 ( .A(n288), .B(n551), .Z(n340) );
  AN2SVTX4 U403 ( .A(n1632), .B(n1617), .Z(n1631) );
  BFSVTX2 U404 ( .A(n1580), .Z(n1778) );
  F_MUX21NSVTX0H U405 ( .A(n1588), .B(n1587), .S(n1069), .Z(n1589) );
  NR2ASVTX4 U406 ( .A(n1620), .B(n1591), .Z(n1626) );
  NR2SVTX6 U407 ( .A(n1591), .B(n1576), .Z(n1577) );
  ND2SVTX4 U408 ( .A(n1749), .B(n1463), .Z(n1501) );
  IVSVTX2 U409 ( .A(n373), .Z(n371) );
  IVSVTX2 U410 ( .A(n369), .Z(n1512) );
  IVSVTX2 U411 ( .A(n1775), .Z(n289) );
  ND2ASVTX6 U412 ( .A(n1566), .B(n738), .Z(n1613) );
  IVSVTX4 U413 ( .A(n530), .Z(n370) );
  NR2SVTX2 U414 ( .A(n1677), .B(n1676), .Z(n1575) );
  AO6SVTX6 U415 ( .A(n1774), .B(n1773), .C(n1217), .Z(n1218) );
  ND2ASVTX4 U416 ( .A(n1547), .B(n1599), .Z(n1612) );
  B_IVSVTX1 U417 ( .A(n1450), .Z(n600) );
  ND2ASVTX6 U418 ( .A(n1258), .B(n1098), .Z(n1440) );
  IVSVTX6 U419 ( .A(n1768), .Z(n1765) );
  ND2ASVTX6 U420 ( .A(n1223), .B(n485), .Z(n1782) );
  ND2ASVTX6 U421 ( .A(n1488), .B(n1487), .Z(n1697) );
  ND3SVTX6 U422 ( .A(n1552), .B(n1551), .C(n1550), .Z(n738) );
  ND2ASVTX4 U423 ( .A(n278), .B(n654), .Z(n599) );
  ND4ABSVTX2 U424 ( .A(n1505), .B(n757), .C(n1421), .D(n1420), .Z(n694) );
  ND4ABSVTX4 U425 ( .A(n1262), .B(n644), .C(n645), .D(n588), .Z(n1769) );
  IVSVTX2 U426 ( .A(n1487), .Z(n1475) );
  IVSVTX0H U427 ( .A(n1220), .Z(n1223) );
  IVSVTX2 U428 ( .A(n589), .Z(n1117) );
  ND2ASVTX6 U429 ( .A(n769), .B(n1489), .Z(n1491) );
  IVSVTX0H U430 ( .A(n1486), .Z(n1488) );
  IVSVTX2 U431 ( .A(n1494), .Z(n1496) );
  B_ND2SVTX2 U432 ( .A(n1203), .B(n1202), .Z(n1204) );
  NR2ASVTX4 U433 ( .A(n1211), .B(n1210), .Z(n1805) );
  ND2SVTX2 U434 ( .A(n1677), .B(n1119), .Z(n1552) );
  ND2SVTX6 U435 ( .A(n541), .B(n540), .Z(n518) );
  IVSVTX2 U436 ( .A(n1650), .Z(n1566) );
  IVSVTX0H U437 ( .A(n1493), .Z(n1494) );
  ND3SVTX2 U438 ( .A(n1186), .B(n1185), .C(n1184), .Z(n1208) );
  IVSVTX0H U439 ( .A(n302), .Z(n1118) );
  IVSVTX2 U440 ( .A(n1451), .Z(n298) );
  ND3ABSVTX6 U441 ( .A(n437), .B(n292), .C(n801), .Z(n1430) );
  IVSVTX0H U442 ( .A(n1258), .Z(n1099) );
  NR2ASVTX1 U443 ( .A(n304), .B(n475), .Z(n1197) );
  IVSVTX0H U444 ( .A(n1199), .Z(n690) );
  IVSVTX2 U445 ( .A(n1143), .Z(n1144) );
  B_IVSVTX1 U446 ( .A(n1222), .Z(n479) );
  ND3SVTX4 U447 ( .A(n662), .B(n661), .C(n663), .Z(n488) );
  IVSVTX2 U448 ( .A(n1425), .Z(n1426) );
  IVSVTX2 U449 ( .A(n279), .Z(n277) );
  AN2SVTX2 U450 ( .A(n1499), .B(n1119), .Z(n769) );
  B_ND2SVTX2 U451 ( .A(n1483), .B(n1213), .Z(n364) );
  ENSVTX6 U452 ( .A(n295), .B(n546), .Z(n654) );
  IVSVTX4 U453 ( .A(n1555), .Z(n717) );
  AO7CSVTX2 U454 ( .A(n294), .B(n1542), .C(n1478), .Z(n669) );
  B_ND2SVTX2 U455 ( .A(n1211), .B(n956), .Z(n662) );
  IVSVTX4 U456 ( .A(n746), .Z(n712) );
  CTBUFSVTX2 U457 ( .A(n660), .Z(n242) );
  AO6SVTX6 U458 ( .A(n1267), .B(n282), .C(n270), .Z(n639) );
  ND3ASVTX4 U459 ( .A(n1094), .B(n1200), .C(n502), .Z(n1196) );
  B_IVSVTX1 U460 ( .A(n776), .Z(n260) );
  ND2ASVTX4 U461 ( .A(n1647), .B(n272), .Z(n642) );
  AO2SVTX4 U462 ( .A(n1212), .B(n282), .C(n302), .D(n1119), .Z(n365) );
  IVSVTX6 U463 ( .A(n1720), .Z(n279) );
  IVSVTX2 U464 ( .A(n502), .Z(n1211) );
  IVSVTX2 U465 ( .A(n1264), .Z(n1142) );
  CTIVSVTX6 U466 ( .A(n1402), .Z(n618) );
  ND3ABSVTX6 U467 ( .A(n1609), .B(n1585), .C(n641), .Z(n481) );
  BFSVTX2 U468 ( .A(n1230), .Z(n302) );
  B_IVSVTX1 U469 ( .A(n1209), .Z(n1201) );
  NR2SVTX4 U470 ( .A(n1451), .B(n1542), .Z(n482) );
  ND2SVTX2 U471 ( .A(n1253), .B(n1252), .Z(n1486) );
  IVSVTX4 U472 ( .A(n745), .Z(n560) );
  IVSVTX4 U473 ( .A(n1259), .Z(n228) );
  ND2ASVTX4 U474 ( .A(n1135), .B(n1119), .Z(n1222) );
  IVSVTX0H U475 ( .A(n1203), .Z(n219) );
  IVSVTX8 U476 ( .A(n1647), .Z(n1402) );
  IVSVTX2 U477 ( .A(n1483), .Z(n745) );
  IVSVTX2 U478 ( .A(n615), .Z(n614) );
  IVSVTX10 U479 ( .A(n1381), .Z(n1555) );
  AN2SVTX6 U480 ( .A(n1162), .B(n1110), .Z(n1159) );
  ND3SVTX6 U481 ( .A(n1470), .B(n1469), .C(n271), .Z(n1471) );
  IVSVTX2 U482 ( .A(n1244), .Z(n296) );
  F_ND2ASVTX2 U483 ( .A(n1179), .B(n1178), .Z(n1209) );
  IVSVTX2 U484 ( .A(n1258), .Z(n217) );
  AO4SVTX2 U485 ( .A(n447), .B(n446), .C(n475), .D(n1189), .Z(n502) );
  MUX21NSVTX2 U486 ( .A(n1068), .B(n1251), .S(n1069), .Z(n1252) );
  ND2ASVTX6 U487 ( .A(n1412), .B(n1415), .Z(n1585) );
  ND3ABSVTX6 U488 ( .A(n1454), .B(n1453), .C(n1452), .Z(n1499) );
  IVSVTX0H U489 ( .A(n1187), .Z(n447) );
  NR2ASVTX1 U490 ( .A(n1520), .B(n1299), .Z(n1528) );
  IVSVTX2 U491 ( .A(n1215), .Z(n300) );
  IVSVTX2 U492 ( .A(n265), .Z(n1155) );
  IVSVTX0H U493 ( .A(n1313), .Z(n1189) );
  IVSVTX6 U494 ( .A(n1647), .Z(n746) );
  IVSVTX0H U495 ( .A(n1245), .Z(n1248) );
  BFSVTX2 U496 ( .A(n1190), .Z(n360) );
  IVSVTX0H U497 ( .A(n1246), .Z(n1247) );
  ENSVTX6 U498 ( .A(n1162), .B(n1256), .Z(n1183) );
  AO7SVTX1 U499 ( .A(n1009), .B(n1176), .C(n1175), .Z(n1179) );
  AN2SVTX2 U500 ( .A(n1521), .B(n257), .Z(n621) );
  IVSVTX4 U501 ( .A(n1429), .Z(n292) );
  NR3ASVTX4 U502 ( .A(n562), .B(n1466), .C(n563), .Z(n1089) );
  IVSVTX0H U503 ( .A(n500), .Z(n235) );
  IVSVTX0H U504 ( .A(n1009), .Z(n304) );
  IVSVTX10 U505 ( .A(n956), .Z(n1647) );
  IVSVTX6 U506 ( .A(n634), .Z(n1429) );
  NR3SVTX6 U507 ( .A(n1115), .B(n1170), .C(n1256), .Z(n1116) );
  OR2SVTX2 U508 ( .A(n1113), .B(n1114), .Z(n1220) );
  AO4SVTX6 U509 ( .A(n454), .B(n1147), .C(n1151), .D(n1152), .Z(n1244) );
  NR2SVTX2 U510 ( .A(n1393), .B(n1392), .Z(n1397) );
  AO4SVTX4 U511 ( .A(n585), .B(O[27]), .C(n285), .D(n1398), .Z(n1410) );
  IVSVTX1 U512 ( .A(n303), .Z(n226) );
  IVSVTX4 U513 ( .A(n633), .Z(n634) );
  NR2SVTX2 U514 ( .A(n389), .B(n1124), .Z(n898) );
  B_ND2SVTX2 U515 ( .A(n500), .B(n602), .Z(n772) );
  ND2SVTX4 U516 ( .A(n1413), .B(n1394), .Z(n637) );
  AO4SVTX4 U517 ( .A(n1312), .B(n1299), .C(n1357), .D(n622), .Z(n1533) );
  IVSVTX4 U518 ( .A(n232), .Z(n1399) );
  ND3ABSVTX4 U519 ( .A(O[28]), .B(n996), .C(n1413), .Z(n1167) );
  BFSVTX4 U520 ( .A(n703), .Z(n556) );
  IVSVTX2 U521 ( .A(n1414), .Z(n602) );
  IVSVTX0H U522 ( .A(n1403), .Z(n1404) );
  ND2ASVTX6 U523 ( .A(n729), .B(n1106), .Z(n1128) );
  CTIVSVTX2 U524 ( .A(n1156), .Z(n1158) );
  IVSVTX0H U525 ( .A(n1165), .Z(n463) );
  AN2SVTX4 U526 ( .A(n1154), .B(n561), .Z(n265) );
  NR3ABSVTX6 U527 ( .A(n1348), .B(n1349), .C(n1347), .Z(n1417) );
  CTBUFSVTX2 U528 ( .A(n648), .Z(n499) );
  ND3SVTX2 U529 ( .A(n1139), .B(n1138), .C(n1525), .Z(n1141) );
  AO4SVTX6 U530 ( .A(n978), .B(n790), .C(n664), .D(n1343), .Z(n1464) );
  BFSVTX4 U531 ( .A(n1365), .Z(n486) );
  ND2ASVTX6 U532 ( .A(n664), .B(n1398), .Z(n1389) );
  ND2ASVTX6 U533 ( .A(n1334), .B(n1371), .Z(n1351) );
  ND2SVTX2 U534 ( .A(n968), .B(n1448), .Z(n978) );
  AO7SVTX2 U535 ( .A(n276), .B(n1291), .C(n1290), .Z(n1300) );
  ND2SVTX6 U536 ( .A(n1321), .B(n1091), .Z(n678) );
  IVSVTX0H U537 ( .A(n1129), .Z(n1130) );
  ND2SVTX2 U538 ( .A(n1123), .B(n1122), .Z(n1126) );
  CTIVSVTX2 U539 ( .A(n357), .Z(n249) );
  IVSVTX2 U540 ( .A(n1140), .Z(n703) );
  CTBUFSVTX4 U541 ( .A(n1043), .Z(n579) );
  IVSVTX2 U542 ( .A(n632), .Z(n325) );
  B_ND2SVTX2 U543 ( .A(n1106), .B(n1105), .Z(n1102) );
  NR3SVTX6 U544 ( .A(n385), .B(n1181), .C(n734), .Z(n508) );
  BFSVTX2 U545 ( .A(n1045), .Z(n241) );
  NR3SVTX4 U546 ( .A(n1446), .B(n1447), .C(n892), .Z(n1453) );
  ND2SVTX2 U547 ( .A(n251), .B(n250), .Z(n713) );
  NR2SVTX4 U548 ( .A(n1411), .B(n1412), .Z(n627) );
  AO2SVTX4 U549 ( .A(n624), .B(n730), .C(n503), .D(n322), .Z(n1531) );
  CTIVSVTX2 U550 ( .A(n962), .Z(n657) );
  IVSVTX2 U551 ( .A(n1140), .Z(n601) );
  ND2SVTX6 U552 ( .A(n800), .B(n1358), .Z(n1414) );
  CTIVSVTX2 U553 ( .A(n779), .Z(n250) );
  ND2SVTX4 U554 ( .A(n1445), .B(n1408), .Z(n1337) );
  NR2SVTX6 U555 ( .A(n1334), .B(n1299), .Z(n632) );
  ND3SVTX4 U556 ( .A(O[29]), .B(n1082), .C(n395), .Z(n483) );
  ND3SVTX6 U557 ( .A(n1085), .B(n305), .C(n1084), .Z(n375) );
  ND3SVTX6 U558 ( .A(n693), .B(n1052), .C(n1111), .Z(n1053) );
  IVSVTX4 U559 ( .A(n624), .Z(n715) );
  F_ND2ASVTX2 U560 ( .A(n985), .B(n1105), .Z(n733) );
  ND2ASVTX6 U561 ( .A(n1074), .B(n1366), .Z(n1148) );
  IVSVTX1 U562 ( .A(n1367), .Z(n1341) );
  ND2ASVTX6 U563 ( .A(n658), .B(n1324), .Z(n1149) );
  IVSVTX6 U564 ( .A(n773), .Z(n305) );
  IVSVTX10 U565 ( .A(n985), .Z(n1525) );
  CTBUFSVTX4 U566 ( .A(n651), .Z(n509) );
  ND3SVTX2 U567 ( .A(n1122), .B(n1123), .C(n957), .Z(n1035) );
  ND3SVTX4 U568 ( .A(n1137), .B(n1070), .C(n1339), .Z(n1245) );
  NR2SVTX2 U569 ( .A(n308), .B(n1044), .Z(n1129) );
  ND3ABSVTX4 U570 ( .A(n1361), .B(n497), .C(n974), .Z(n1403) );
  AO7SVTX2 U571 ( .A(n1012), .B(n903), .C(n1275), .Z(n1315) );
  BFSVTX2 U572 ( .A(n1033), .Z(n212) );
  AO3SVTX6 U573 ( .A(n1042), .B(n1041), .C(n1049), .D(n1048), .Z(n693) );
  F_IVSVTX1 U574 ( .A(n895), .Z(n896) );
  IVSVTX6 U575 ( .A(n1339), .Z(n1447) );
  IVSVTX2 U576 ( .A(n1137), .Z(n1074) );
  IVSVTX4 U577 ( .A(O[29]), .Z(n307) );
  IVSVTX2 U578 ( .A(n1274), .Z(n1275) );
  IVSVTX4 U579 ( .A(n452), .Z(n1313) );
  ND2SVTX2 U580 ( .A(n1059), .B(n1058), .Z(n1076) );
  ND3ASVTX6 U581 ( .A(n1283), .B(n1282), .C(n1281), .Z(n1360) );
  IVSVTX8 U582 ( .A(n229), .Z(n624) );
  ND3SVTX4 U583 ( .A(n895), .B(n1051), .C(n1050), .Z(n1104) );
  AO4SVTX4 U584 ( .A(n582), .B(n1044), .C(n1043), .D(n1045), .Z(n583) );
  AO6SVTX4 U585 ( .A(n724), .B(n882), .C(n759), .Z(n907) );
  IVSVTX2 U586 ( .A(n1043), .Z(n582) );
  AO7SVTX4 U587 ( .A(n498), .B(n497), .C(n1028), .Z(n501) );
  ND3ABSVTX4 U588 ( .A(n1031), .B(O[31]), .C(n1325), .Z(n231) );
  ND2SVTX2 U589 ( .A(n990), .B(n992), .Z(n892) );
  IVSVTX4 U590 ( .A(n1044), .Z(n514) );
  NR2ASVTX4 U591 ( .A(n933), .B(n586), .Z(n1274) );
  ND2SVTX2 U592 ( .A(n1325), .B(n971), .Z(n973) );
  IVSVTX4 U593 ( .A(n949), .Z(n308) );
  ND2SVTX4 U594 ( .A(n1013), .B(n1043), .Z(n652) );
  NR2ASVTX1 U595 ( .A(n1277), .B(n587), .Z(n1283) );
  F_ND2ASVTX2 U596 ( .A(n964), .B(n673), .Z(n966) );
  AO4SVTX4 U597 ( .A(n497), .B(n997), .C(n996), .D(n306), .Z(n685) );
  AO7SVTX6 U598 ( .A(n912), .B(O[31]), .C(n650), .Z(n913) );
  AO2SVTX4 U599 ( .A(n606), .B(n605), .C(n777), .D(n940), .Z(n608) );
  MUX21NSVTX6 U600 ( .A(n1006), .B(N[0]), .S(n1019), .Z(n1188) );
  ND2SVTX2 U601 ( .A(n923), .B(n1292), .Z(n319) );
  ND2ASVTX1 U602 ( .A(n276), .B(n1294), .Z(n1180) );
  IVSVTX10 U603 ( .A(n722), .Z(O[29]) );
  IVSVTX1 U604 ( .A(n852), .Z(n691) );
  AO6ABSVTX6 U605 ( .A(n980), .B(n424), .C(n979), .Z(n997) );
  BFSVTX8 U606 ( .A(n1072), .Z(n327) );
  IVSVTX0H U607 ( .A(n311), .Z(n334) );
  IVSVTX0H U608 ( .A(n1279), .Z(n1280) );
  ND3ASVTX2 U609 ( .A(n812), .B(n587), .C(n752), .Z(n1064) );
  ND3SVTX4 U610 ( .A(n1059), .B(n1123), .C(n1058), .Z(n1050) );
  IVSVTX4 U611 ( .A(n306), .Z(n417) );
  NR2SVTX1 U612 ( .A(n1031), .B(n1030), .Z(n1032) );
  ND3ABSVTX4 U613 ( .A(n872), .B(n243), .C(O[31]), .Z(n1332) );
  IVSVTX0H U614 ( .A(n927), .Z(n970) );
  NR3ABSVTX6 U615 ( .A(n1003), .B(n754), .C(n1176), .Z(n441) );
  BFSVTX0H U616 ( .A(N[15]), .Z(n933) );
  BFSVTX0H U617 ( .A(N[16]), .Z(n959) );
  ND2ASVTX6 U618 ( .A(n1279), .B(n932), .Z(n1047) );
  ND2ASVTX6 U619 ( .A(n812), .B(n426), .Z(n1123) );
  BFSVTX0H U620 ( .A(n680), .Z(n679) );
  IVSVTX2 U621 ( .A(n754), .Z(n423) );
  AN2SVTX6 U622 ( .A(n516), .B(n894), .Z(n418) );
  ND2SVTX4 U623 ( .A(n1021), .B(n462), .Z(n1025) );
  IVSVTX0H U624 ( .A(n922), .Z(n923) );
  IVSVTX10 U625 ( .A(n737), .Z(n948) );
  ND2ASVTX4 U626 ( .A(n1293), .B(n958), .Z(n1061) );
  ND3ABSVTX4 U627 ( .A(n1279), .B(n984), .C(n656), .Z(n1176) );
  BFSVTX0H U628 ( .A(N[13]), .Z(n1284) );
  IVSVTX0H U629 ( .A(n1020), .Z(n243) );
  CTIVSVTX4 U630 ( .A(n947), .Z(n591) );
  IVSVTX4 U631 ( .A(n425), .Z(n424) );
  NR2ASVTX4 U632 ( .A(N[4]), .B(n1285), .Z(n396) );
  NR2ASVTX6 U633 ( .A(n1038), .B(n1037), .Z(n1083) );
  CTIVSVTX2 U634 ( .A(N[3]), .Z(n1279) );
  ND2ASVTX4 U635 ( .A(n1293), .B(n1292), .Z(n1328) );
  ND3SVTX6 U636 ( .A(N[1]), .B(n587), .C(n752), .Z(n775) );
  ND4SVTX4 U637 ( .A(n943), .B(n1017), .C(n944), .D(n535), .Z(n317) );
  IVSVTX6 U638 ( .A(n725), .Z(n945) );
  IVSVTX6 U639 ( .A(n910), .Z(n911) );
  IVSVTX6 U640 ( .A(n983), .Z(n894) );
  IVSVTX1 U641 ( .A(N[12]), .Z(n1293) );
  IVSVTX2 U642 ( .A(N[0]), .Z(n276) );
  ND3SVTX6 U643 ( .A(n981), .B(n484), .C(n1017), .Z(n982) );
  ND3ASVTX4 U644 ( .A(n1012), .B(n958), .C(n470), .Z(n469) );
  BFSVTX2 U645 ( .A(N[4]), .Z(n1326) );
  CTIVSVTX2 U646 ( .A(N[1]), .Z(n1005) );
  BFSVTX4 U647 ( .A(n1018), .Z(n515) );
  IVSVTX2 U648 ( .A(n1017), .Z(n470) );
  IVSVTX10 U649 ( .A(n587), .Z(n1294) );
  IVSVTX2 U650 ( .A(n1038), .Z(n1012) );
  ND3SVTX6 U651 ( .A(n990), .B(n991), .C(n992), .Z(n1075) );
  IVSVTX0H U652 ( .A(n1278), .Z(n888) );
  NR2SVTX2 U653 ( .A(n675), .B(n870), .Z(n505) );
  BFSVTX2 U654 ( .A(N[2]), .Z(n981) );
  IVSVTX6 U655 ( .A(n872), .Z(n310) );
  BFSVTX4 U656 ( .A(n868), .Z(n484) );
  NR2SVTX6 U657 ( .A(n831), .B(n830), .Z(n909) );
  BFSVTX2 U658 ( .A(N[7]), .Z(n1038) );
  ND3ABSVTX6 U659 ( .A(n845), .B(n869), .C(n857), .Z(n831) );
  IVSVTX2 U660 ( .A(n812), .Z(n720) );
  F_ND2ASVTX2 U661 ( .A(n672), .B(n880), .Z(n884) );
  ND4SVTX2 U662 ( .A(N[1]), .B(n1031), .C(n827), .D(n828), .Z(n811) );
  BFSVTX6 U663 ( .A(N[5]), .Z(n1020) );
  IVSVTX6 U664 ( .A(n448), .Z(n860) );
  NR2SVTX4 U665 ( .A(n841), .B(n842), .Z(n850) );
  NR2ASVTX4 U666 ( .A(N[3]), .B(n675), .Z(n829) );
  CTIVSVTX2 U667 ( .A(n825), .Z(n826) );
  NR2SVTX6 U668 ( .A(n818), .B(n868), .Z(n547) );
  B_ND2SVTX2 U669 ( .A(n902), .B(n760), .Z(n820) );
  ND3SVTX6 U670 ( .A(n901), .B(n312), .C(n1018), .Z(n865) );
  IVSVTX2 U671 ( .A(N[6]), .Z(n812) );
  IVSVTX2 U672 ( .A(n870), .Z(n761) );
  NR2SVTX4 U673 ( .A(N[12]), .B(N[13]), .Z(n881) );
  IVSVTX8 U674 ( .A(n849), .Z(n368) );
  IVSVTX6 U675 ( .A(n809), .Z(n880) );
  IVSVTX2 U676 ( .A(n862), .Z(n864) );
  NR2SVTX6 U677 ( .A(n675), .B(n845), .Z(n847) );
  CTBUFSVTX4 U678 ( .A(n863), .Z(n321) );
  IVSVTX2 U679 ( .A(n902), .Z(n704) );
  IVSVTX1 U680 ( .A(N[31]), .Z(n840) );
  NR2SVTX4 U681 ( .A(N[25]), .B(N[27]), .Z(n549) );
  NR2SVTX4 U682 ( .A(N[18]), .B(N[30]), .Z(n804) );
  NR2SVTX6 U683 ( .A(N[31]), .B(N[28]), .Z(n655) );
  IVSVTX6 U684 ( .A(N[28]), .Z(n680) );
  IVSVTX10 U685 ( .A(N[29]), .Z(n924) );
  IVSVTX8 U686 ( .A(n211), .Z(n214) );
  AO7SVTX8 U687 ( .A(n1385), .B(n1384), .C(n1383), .Z(n211) );
  NR2SVTX4 U688 ( .A(n1238), .B(n1714), .Z(n1436) );
  ND2SVTX4 U689 ( .A(n1790), .B(n1797), .Z(n1714) );
  AO7SVTX4 U690 ( .A(n1291), .B(n917), .C(n259), .Z(n918) );
  IVSVTX6 U691 ( .A(n1727), .Z(n1684) );
  AO7SVTX8 U692 ( .A(n1739), .B(n531), .C(n1670), .Z(n1727) );
  AO5SVTX6 U693 ( .A(n1637), .B(n1638), .C(n378), .Z(n1618) );
  IVSVTX12 U694 ( .A(n1646), .Z(n764) );
  ND3ASVTX8 U695 ( .A(n1574), .B(n764), .C(n401), .Z(n393) );
  IVSVTX8 U696 ( .A(n261), .Z(n1664) );
  ENSVTX6 U697 ( .A(n1228), .B(n1116), .Z(n1120) );
  ND2SVTX6 U698 ( .A(n399), .B(n400), .Z(n1673) );
  ND3ABSVTX8 U699 ( .A(n1255), .B(n1256), .C(n1089), .Z(n1090) );
  ENSVTX8 U700 ( .A(n1220), .B(n366), .Z(n1213) );
  ND3SVTX8 U701 ( .A(n424), .B(n775), .C(n710), .Z(n1024) );
  AO7SVTX6 U702 ( .A(n579), .B(n581), .C(n580), .Z(n1107) );
  IVSVTX6 U703 ( .A(n1124), .Z(n256) );
  BFSVTX1 U704 ( .A(n457), .Z(n213) );
  ND3ASVTX6 U705 ( .A(n722), .B(n1370), .C(n1124), .Z(n891) );
  AO7SVTX8 U706 ( .A(n712), .B(n233), .C(n214), .Z(n1630) );
  IVSVTX12 U707 ( .A(n777), .Z(n1325) );
  ND2SVTX4 U708 ( .A(n985), .B(n501), .Z(n1029) );
  AO4SVTX8 U709 ( .A(n407), .B(n408), .C(n406), .D(n1526), .Z(n951) );
  IVSVTX4 U710 ( .A(n1254), .Z(n216) );
  ND3SVTX6 U711 ( .A(n217), .B(n216), .C(n512), .Z(n1257) );
  AO7ABSVTX6 U712 ( .A(n541), .B(n1477), .C(n1474), .Z(n1487) );
  ND3SVTX8 U713 ( .A(n424), .B(n1014), .C(n1015), .Z(n1027) );
  F_ND2ASVTX2 U714 ( .A(n912), .B(n872), .Z(n1014) );
  BFSVTX1 U715 ( .A(n1435), .Z(n218) );
  OR2SVTX4 U716 ( .A(n219), .B(n709), .Z(n661) );
  AO7ABSVTX4 U717 ( .A(n220), .B(n1574), .C(n221), .Z(n392) );
  IVSVTX4 U718 ( .A(n1119), .Z(n1808) );
  AO5SVTX6 U719 ( .A(n1655), .B(n224), .C(n1654), .Z(n261) );
  ND4ASVTX8 U720 ( .A(n330), .B(n848), .C(n847), .D(n846), .Z(n459) );
  IVSVTX4 U721 ( .A(n236), .Z(n275) );
  IVSVTX10 U722 ( .A(n818), .Z(n312) );
  ENSVTX8 U723 ( .A(n780), .B(n222), .Z(O[23]) );
  AO6SVTX4 U724 ( .A(n1741), .B(n286), .C(n223), .Z(n222) );
  IVSVTX10 U725 ( .A(n681), .Z(n576) );
  IVSVTX10 U726 ( .A(n1109), .Z(n1110) );
  ND3ABSVTX6 U727 ( .A(n276), .B(O[31]), .C(n674), .Z(n522) );
  AO6CSVTX8 U728 ( .A(n1249), .B(n1250), .C(n1140), .Z(n1088) );
  IVSVTX6 U729 ( .A(n1574), .Z(n1718) );
  IVSVTX6 U730 ( .A(n565), .Z(n322) );
  ND2SVTX4 U731 ( .A(n226), .B(n225), .Z(n1380) );
  NR2SVTX4 U732 ( .A(n585), .B(n1414), .Z(n225) );
  AO7SVTX8 U733 ( .A(n712), .B(n1269), .C(n227), .Z(n676) );
  AO6SVTX8 U734 ( .A(n578), .B(n282), .C(n228), .Z(n227) );
  AO7SVTX4 U735 ( .A(n1492), .B(n1697), .C(n1690), .Z(n337) );
  NR2SVTX4 U736 ( .A(n1490), .B(n1484), .Z(n1492) );
  ND3ABSVTX8 U737 ( .A(N[27]), .B(N[25]), .C(n414), .Z(n822) );
  CTIVSVTX4 U738 ( .A(n1455), .Z(n1468) );
  ND3ASVTX8 U739 ( .A(n1574), .B(n1628), .C(n764), .Z(n255) );
  IVSVTX12 U740 ( .A(n1356), .Z(n1522) );
  CTIVSVTX4 U741 ( .A(n388), .Z(n513) );
  IVSVTX4 U742 ( .A(n1366), .Z(n229) );
  NR2ASVTX2 U743 ( .A(n1003), .B(n737), .Z(n987) );
  IVSVTX4 U744 ( .A(n1574), .Z(n383) );
  AO7SVTX8 U745 ( .A(n657), .B(n715), .C(n1330), .Z(n1331) );
  AO7ABSVTX6 U746 ( .A(n1300), .B(n322), .C(n1298), .Z(n1394) );
  ENSVTX8 U747 ( .A(n296), .B(n1153), .Z(n573) );
  AO7SVTX6 U748 ( .A(n864), .B(n321), .C(n705), .Z(n866) );
  ND3SVTX8 U749 ( .A(n680), .B(n650), .C(n316), .Z(n836) );
  NR2ASVTX8 U750 ( .A(n968), .B(n1343), .Z(n1344) );
  ND2SVTX6 U751 ( .A(n1531), .B(n1529), .Z(n1396) );
  ND2ASVTX8 U752 ( .A(n1647), .B(n1120), .Z(n686) );
  ND3SVTX8 U753 ( .A(n1200), .B(n283), .C(n1617), .Z(n1186) );
  ND3SVTX8 U754 ( .A(n967), .B(n966), .C(n231), .Z(n1367) );
  ND3SVTX8 U755 ( .A(n483), .B(n891), .C(n890), .Z(n1251) );
  ND3SVTX6 U756 ( .A(n1390), .B(n1389), .C(n706), .Z(n232) );
  ENSVTX6 U757 ( .A(n1677), .B(n1382), .Z(n233) );
  IVSVTX4 U758 ( .A(n1409), .Z(n428) );
  ND2SVTX4 U759 ( .A(n1480), .B(n1481), .Z(n1482) );
  ND3SVTX6 U760 ( .A(n341), .B(n342), .C(n1459), .Z(n1480) );
  ND2SVTX4 U761 ( .A(n332), .B(n1198), .Z(n734) );
  IVSVTX12 U762 ( .A(n234), .Z(n1285) );
  ND3SVTX8 U763 ( .A(n807), .B(n806), .C(n805), .Z(n234) );
  IVSVTX10 U764 ( .A(n822), .Z(n1018) );
  NR3SVTX8 U765 ( .A(n1109), .B(n1255), .C(n1254), .Z(n1243) );
  ND3SVTX6 U766 ( .A(n1244), .B(n1242), .C(n1241), .Z(n1254) );
  F_ND2ASVTX2 U767 ( .A(n235), .B(n1532), .Z(n1310) );
  ND2ASVTX8 U768 ( .A(n1317), .B(n486), .Z(n1307) );
  AO4SVTX4 U769 ( .A(n1718), .B(n1119), .C(n753), .D(n1646), .Z(n236) );
  ND3SVTX8 U770 ( .A(n1150), .B(n1245), .C(n1148), .Z(n1079) );
  IVSVTX4 U771 ( .A(n237), .Z(n785) );
  ND3ASVTX6 U772 ( .A(n1388), .B(n297), .C(n1377), .Z(n237) );
  ND3ABSVTX8 U773 ( .A(n945), .B(n317), .C(n591), .Z(n592) );
  ND2SVTX4 U774 ( .A(n1273), .B(n325), .Z(n1376) );
  IVSVTX6 U775 ( .A(n748), .Z(n1299) );
  IVSVTX4 U776 ( .A(n239), .Z(n1590) );
  ND2SVTX4 U777 ( .A(n1521), .B(n748), .Z(n239) );
  AN2SVTX8 U778 ( .A(n1339), .B(n1387), .Z(n748) );
  ND2SVTX4 U779 ( .A(n240), .B(n765), .Z(n384) );
  AN2SVTX4 U780 ( .A(n294), .B(n1513), .Z(n801) );
  ND3SVTX8 U781 ( .A(n395), .B(n664), .C(n471), .Z(n666) );
  ND2ASVTX8 U782 ( .A(n1647), .B(n1473), .Z(n640) );
  AO3SVTX8 U783 ( .A(n1269), .B(n278), .C(n1268), .D(n796), .Z(n388) );
  ND2ASVTX8 U784 ( .A(n1238), .B(n1712), .Z(n1240) );
  IVSVTX8 U785 ( .A(n255), .Z(n1656) );
  ND2ASVTX8 U786 ( .A(n1106), .B(n244), .Z(n344) );
  IVSVTX4 U787 ( .A(n1526), .Z(n244) );
  AO6SVTX6 U788 ( .A(n1292), .B(n959), .C(n913), .Z(n1290) );
  BFSVTX1 U789 ( .A(n1745), .Z(n245) );
  NR2SVTX4 U790 ( .A(n246), .B(n577), .Z(n259) );
  AO7SVTX6 U791 ( .A(n1293), .B(O[31]), .C(n679), .Z(n246) );
  AO6SVTX2 U792 ( .A(n1517), .B(n1625), .C(n1516), .Z(n1518) );
  AO7SVTX6 U793 ( .A(n248), .B(n247), .C(n1160), .Z(n338) );
  IVSVTX4 U794 ( .A(n788), .Z(n247) );
  ND2SVTX4 U795 ( .A(n358), .B(n249), .Z(n248) );
  IVSVTX6 U796 ( .A(n1424), .Z(n633) );
  ND3SVTX8 U797 ( .A(n627), .B(n628), .C(n626), .Z(n1424) );
  IVSVTX4 U798 ( .A(n565), .Z(n251) );
  AO6SVTX6 U799 ( .A(n1062), .B(n1061), .C(n327), .Z(n1066) );
  ND2SVTX4 U800 ( .A(n253), .B(n471), .Z(n800) );
  IVSVTX4 U801 ( .A(n1357), .Z(n253) );
  ND3SVTX6 U802 ( .A(n254), .B(n520), .C(n871), .Z(n885) );
  NR2SVTX4 U803 ( .A(n675), .B(n869), .Z(n254) );
  AO7SVTX8 U804 ( .A(n1610), .B(n1613), .C(n1612), .Z(n1622) );
  ND3SVTX6 U805 ( .A(n1085), .B(n1081), .C(n1084), .Z(n1152) );
  ND2SVTX4 U806 ( .A(n256), .B(n376), .Z(n1081) );
  ND4SVTX4 U807 ( .A(n1546), .B(n1547), .C(n1555), .D(n641), .Z(n1548) );
  IVSVTX4 U808 ( .A(n676), .Z(n1261) );
  AO7SVTX6 U809 ( .A(n1490), .B(n1491), .C(n411), .Z(n1690) );
  ND3SVTX8 U810 ( .A(n1097), .B(n766), .C(n338), .Z(n709) );
  ND2ASVTX8 U811 ( .A(n950), .B(n575), .Z(n766) );
  ND2SVTX6 U812 ( .A(n1367), .B(n471), .Z(n1448) );
  AO7SVTX6 U813 ( .A(n570), .B(n596), .C(n285), .Z(n595) );
  IVSVTX4 U814 ( .A(n1499), .Z(n1472) );
  IVSVTX6 U815 ( .A(n287), .Z(n432) );
  ND2SVTX8 U816 ( .A(n1321), .B(n1091), .Z(n1109) );
  ND2SVTX6 U817 ( .A(n1617), .B(n287), .Z(n379) );
  NR2SVTX6 U818 ( .A(N[16]), .B(N[26]), .Z(n316) );
  ND3SVTX8 U819 ( .A(n383), .B(n1634), .C(n1633), .Z(n1654) );
  IVSVTX6 U820 ( .A(n1019), .Z(n743) );
  ENSVTX8 U821 ( .A(n1674), .B(n1673), .Z(n445) );
  BFSVTX6 U822 ( .A(n1371), .Z(n257) );
  AO21SVTX8 U823 ( .A(n615), .B(n613), .C(n610), .D(n1650), .Z(n609) );
  ND4ABSVTX8 U824 ( .A(n1251), .B(n1088), .C(n1086), .D(n1087), .Z(n1466) );
  ND2SVTX4 U825 ( .A(n1679), .B(n258), .Z(n457) );
  ND2ASVTX8 U826 ( .A(n524), .B(n340), .Z(n1583) );
  AO7ABSVTX6 U827 ( .A(n295), .B(n1584), .C(n1583), .Z(n339) );
  AO7ASVTX8 U828 ( .A(n369), .B(n1511), .C(n1510), .Z(n1565) );
  IVSVTX6 U829 ( .A(n1580), .Z(n1506) );
  AO7SVTX8 U830 ( .A(n604), .B(n603), .C(n405), .Z(n1580) );
  AO17SVTX8 U831 ( .A(n429), .B(n430), .C(n381), .D(n1746), .Z(n1642) );
  ND3ASVTX6 U832 ( .A(n260), .B(n645), .C(n588), .Z(n1263) );
  AO6SVTX8 U833 ( .A(n1187), .B(n1276), .C(n1004), .Z(n1008) );
  EO3SVTX8 U834 ( .A(n1655), .B(n1656), .C(n1654), .Z(n1640) );
  IVSVTX4 U835 ( .A(n263), .Z(n270) );
  ND2SVTX4 U836 ( .A(n1119), .B(n1476), .Z(n263) );
  AO7SVTX6 U837 ( .A(n1009), .B(n1188), .C(n1199), .Z(n494) );
  IVSVTX2 U838 ( .A(n441), .Z(n451) );
  ND2SVTX2 U839 ( .A(O[27]), .B(n285), .Z(n636) );
  IVSVTX0H U840 ( .A(n1326), .Z(n1296) );
  ND2SVTX2 U841 ( .A(n1523), .B(n950), .Z(n407) );
  NR2SVTX2 U842 ( .A(n1129), .B(n1140), .Z(n1055) );
  IVSVTX0H U843 ( .A(n972), .Z(n929) );
  IVSVTX2 U844 ( .A(n1620), .Z(n1621) );
  IVSVTX0H U845 ( .A(n941), .Z(n605) );
  AO7ASVTX6 U846 ( .A(n713), .B(n1331), .C(n1413), .Z(n1349) );
  NR2SVTX2 U847 ( .A(n330), .B(n870), .Z(n871) );
  IVSVTX0H U848 ( .A(n1778), .Z(n524) );
  BFSVTX1 U849 ( .A(n1630), .Z(n453) );
  ND3ABSVTX4 U850 ( .A(n1631), .B(n1574), .C(n764), .Z(n399) );
  AO6SVTX1 U851 ( .A(n1784), .B(n1711), .C(n1783), .Z(n1785) );
  F_ND2SVTX0H U852 ( .A(n1755), .B(n1757), .Z(n1760) );
  ENSVTX0H U853 ( .A(n1807), .B(n1806), .Z(O[0]) );
  EOSVTX0H U854 ( .A(n1710), .B(n1709), .Z(O[2]) );
  IVSVTX0H U855 ( .A(n940), .Z(n942) );
  IVSVTX12 U856 ( .A(n853), .Z(n1017) );
  ND2SVTX2 U857 ( .A(n972), .B(n1329), .Z(n264) );
  IVSVTX10 U858 ( .A(n418), .Z(n895) );
  IVSVTX12 U859 ( .A(n1387), .Z(n1140) );
  IVSVTX8 U860 ( .A(n327), .Z(n1000) );
  AN3SVTX4 U861 ( .A(n1128), .B(n500), .C(n1127), .Z(n266) );
  AO17NSVTX8 U862 ( .A(n1137), .B(n1366), .C(n773), .D(n664), .Z(n267) );
  IVSVTX12 U863 ( .A(n387), .Z(n1082) );
  IVSVTX2 U864 ( .A(n1273), .Z(n631) );
  ND2SVTX2 U865 ( .A(n1367), .B(n1371), .Z(n1273) );
  IVSVTX10 U866 ( .A(n620), .Z(n1371) );
  IVSVTX8 U867 ( .A(n1647), .Z(n1483) );
  ND2SVTX2 U868 ( .A(n1585), .B(n1119), .Z(n1450) );
  IVSVTX8 U869 ( .A(n1652), .Z(n294) );
  AO7NSVTX4 U870 ( .A(n1555), .B(n1546), .C(n282), .Z(n268) );
  NR3SVTX2 U871 ( .A(n1468), .B(n1467), .C(n1466), .Z(n271) );
  F_EOSVTX2 U872 ( .A(n284), .B(n1159), .Z(n272) );
  IVSVTX6 U873 ( .A(n1113), .Z(n315) );
  AN2SVTX4 U874 ( .A(n1749), .B(n1463), .Z(n273) );
  IVSVTX8 U875 ( .A(n1542), .Z(n437) );
  F_ENSVTX2 U876 ( .A(n1595), .B(n1594), .Z(n274) );
  ND2SVTX4 U877 ( .A(n768), .B(n394), .Z(n1724) );
  MUX21NSVTX8 U878 ( .A(n413), .B(n412), .S(n1019), .Z(n1187) );
  ND2SVTX2 U879 ( .A(n1525), .B(n1100), .Z(n1101) );
  ND3ABSVTX6 U880 ( .A(n1180), .B(n1070), .C(n1365), .Z(n1198) );
  ND2ASVTX4 U881 ( .A(n1600), .B(n1673), .Z(n398) );
  EOSVTX2 U882 ( .A(n1799), .B(n1798), .Z(O[4]) );
  ND2SVTX4 U883 ( .A(n1509), .B(n1508), .Z(n1608) );
  IVSVTX8 U884 ( .A(n291), .Z(n753) );
  ND2SVTX4 U885 ( .A(n299), .B(n1460), .Z(n1505) );
  CTIVSVTX2 U886 ( .A(n304), .Z(n446) );
  IVSVTX2 U887 ( .A(n968), .Z(n570) );
  IVSVTX8 U888 ( .A(n950), .Z(O[27]) );
  B_ND2SVTX2 U889 ( .A(n1000), .B(n390), .Z(n389) );
  IVSVTX4 U890 ( .A(n1166), .Z(n996) );
  IVSVTX2 U891 ( .A(n854), .Z(n855) );
  B_ND2SVTX2 U892 ( .A(n972), .B(n964), .Z(n814) );
  B_ND2SVTX2 U893 ( .A(n1670), .B(n1663), .Z(n1672) );
  ND2SVTX2 U894 ( .A(n1810), .B(n1809), .Z(n1811) );
  NR2SVTX6 U895 ( .A(n274), .B(n432), .Z(n1596) );
  HA1SVTX6 U896 ( .A(n1609), .B(n1608), .CO(n1629), .S(n1636) );
  ND3ABSVTX6 U897 ( .A(n298), .B(n1507), .C(n695), .Z(n369) );
  ND2ASVTX6 U898 ( .A(n1216), .B(n1214), .Z(n1773) );
  OR2ABSVTX4 U899 ( .A(n712), .B(n293), .Z(n1648) );
  IVSVTX2 U900 ( .A(n1459), .Z(n405) );
  IVSVTX4 U901 ( .A(n1505), .Z(n1459) );
  IVSVTX10 U902 ( .A(n278), .Z(n291) );
  IVSVTX8 U903 ( .A(n282), .Z(n278) );
  ND3SVTX4 U904 ( .A(n1200), .B(n348), .C(n1094), .Z(n362) );
  IVSVTX2 U905 ( .A(n1155), .Z(n348) );
  IVSVTX8 U906 ( .A(n1603), .Z(n1547) );
  ND3ABSVTX6 U907 ( .A(n1169), .B(n1168), .C(n1167), .Z(n1215) );
  ND2SVTX8 U908 ( .A(n939), .B(n1160), .Z(n1190) );
  CTIVSVTX2 U909 ( .A(n1468), .Z(n562) );
  CTIVSVTX2 U910 ( .A(n472), .Z(n566) );
  IVSVTX2 U911 ( .A(n601), .Z(n357) );
  NR2SVTX2 U912 ( .A(O[29]), .B(n877), .Z(n377) );
  ND3SVTX4 U913 ( .A(n1288), .B(n1287), .C(n1286), .Z(n1520) );
  ND2SVTX2 U914 ( .A(n1277), .B(n673), .Z(n935) );
  ND2ASVTX4 U915 ( .A(n861), .B(n1292), .Z(n908) );
  CTIVSVTX4 U916 ( .A(n1291), .Z(n696) );
  IVSVTX10 U917 ( .A(n547), .Z(n872) );
  ND2ASVTX4 U918 ( .A(N[15]), .B(n844), .Z(n848) );
  NR2SVTX6 U919 ( .A(N[20]), .B(N[21]), .Z(n1030) );
  ND2SVTX6 U920 ( .A(n1572), .B(n551), .Z(n1573) );
  FA1SVTX2 U921 ( .A(n453), .B(n1652), .CI(n1651), .CO(n1658), .Z(n1655) );
  ND2SVTX2 U922 ( .A(n1386), .B(n1561), .Z(n1519) );
  ND2SVTX4 U923 ( .A(n1480), .B(n1461), .Z(n552) );
  ND3SVTX6 U924 ( .A(n1549), .B(n268), .C(n1548), .Z(n1550) );
  CTAN2BSVTX4 U925 ( .A(n1652), .B(n709), .Z(n1425) );
  ND2SVTX6 U926 ( .A(n282), .B(n1213), .Z(n687) );
  IVSVTX4 U927 ( .A(n1631), .Z(n293) );
  IVSVTX2 U928 ( .A(n787), .Z(n299) );
  F_ND2ASVTX2 U929 ( .A(n1404), .B(n566), .Z(n787) );
  IVSVTX4 U930 ( .A(n1351), .Z(n303) );
  ND4SVTX6 U931 ( .A(n542), .B(n770), .C(n1289), .D(n324), .Z(n1388) );
  IVSVTX2 U932 ( .A(n416), .Z(n1335) );
  IVSVTX8 U933 ( .A(O[27]), .Z(n285) );
  ND2SVTX4 U934 ( .A(n308), .B(n397), .Z(n492) );
  AO3SVTX6 U935 ( .A(n1291), .B(n1031), .C(n908), .D(n907), .Z(n1523) );
  ND2ASVTX6 U936 ( .A(n989), .B(n988), .Z(n1166) );
  NR2ASVTX4 U937 ( .A(n1020), .B(n1291), .Z(n697) );
  AO7NSVTX4 U938 ( .A(n1296), .B(n903), .C(n1327), .Z(n791) );
  ND2ASVTX4 U939 ( .A(n929), .B(n958), .Z(n710) );
  NR2SVTX6 U940 ( .A(N[14]), .B(N[12]), .Z(n808) );
  BFSVTX6 U941 ( .A(N[19]), .Z(n1277) );
  B_ND2SVTX2 U942 ( .A(n1723), .B(n1682), .Z(n1688) );
  AO7ABSVTX2 U943 ( .A(n1719), .B(n1720), .C(n455), .Z(n1721) );
  ND2SVTX4 U944 ( .A(n1679), .B(n1605), .Z(n1661) );
  EOSVTX2 U945 ( .A(n1760), .B(n1759), .Z(O[14]) );
  B_ND2SVTX2 U946 ( .A(n1659), .B(n1658), .Z(n534) );
  B_ND2SVTX1 U947 ( .A(n751), .B(n1711), .Z(n1715) );
  B_ND2SVTX2 U948 ( .A(n347), .B(n1787), .Z(n1789) );
  ND2ASVTX4 U949 ( .A(n1486), .B(n1475), .Z(n1698) );
  ND2ASVTX4 U950 ( .A(n1235), .B(n1117), .Z(n1797) );
  ND2ASVTX4 U951 ( .A(n1118), .B(n1234), .Z(n1791) );
  ENSVTX4 U952 ( .A(n298), .B(n555), .Z(n554) );
  ND3ABSVTX4 U953 ( .A(n769), .B(n411), .C(n1489), .Z(n1484) );
  ND2ASVTX4 U954 ( .A(n1220), .B(n1222), .Z(n1143) );
  NR2ASVTX4 U955 ( .A(n301), .B(n1202), .Z(n1205) );
  IVSVTX2 U956 ( .A(n1225), .Z(n574) );
  NR2SVTX4 U957 ( .A(n784), .B(n750), .Z(n341) );
  IVSVTX4 U958 ( .A(n1547), .Z(n619) );
  F_ND2ASVTX2 U959 ( .A(n1590), .B(n1589), .Z(n1632) );
  IVSVTX12 U960 ( .A(n1478), .Z(n282) );
  ND3ABSVTX8 U961 ( .A(n1528), .B(n621), .C(n1527), .Z(n1720) );
  IVSVTX4 U962 ( .A(n300), .Z(n283) );
  ND3SVTX4 U963 ( .A(n1149), .B(n1146), .C(n1148), .Z(n454) );
  MUX21NSVTX4 U964 ( .A(n1532), .B(n1587), .S(n500), .Z(n1527) );
  IVSVTX4 U965 ( .A(n1235), .Z(n284) );
  IVSVTX4 U966 ( .A(n733), .Z(n1114) );
  CTIVSVTX4 U967 ( .A(n494), .Z(n386) );
  IVSVTX2 U968 ( .A(n749), .Z(n332) );
  IVSVTX8 U969 ( .A(n410), .Z(n1324) );
  IVSVTX2 U970 ( .A(n1316), .Z(n730) );
  IVSVTX4 U971 ( .A(n950), .Z(n1413) );
  IVSVTX2 U972 ( .A(n503), .Z(n1317) );
  IVSVTX2 U973 ( .A(n1360), .Z(n1312) );
  ND2ASVTX4 U974 ( .A(n692), .B(n691), .Z(n1199) );
  AO7SVTX6 U975 ( .A(n674), .B(n1047), .C(n1046), .Z(n420) );
  ND2ASVTX6 U976 ( .A(n722), .B(n921), .Z(n410) );
  IVSVTX2 U977 ( .A(n1370), .Z(n1336) );
  ND2ASVTX6 U978 ( .A(n1005), .B(n696), .Z(n1306) );
  AO7SVTX6 U979 ( .A(n812), .B(n903), .C(n608), .Z(n1521) );
  IVSVTX4 U980 ( .A(n1039), .Z(n309) );
  AO6CSVTX6 U981 ( .A(n1292), .B(n1032), .C(n793), .Z(n1122) );
  B_ND2SVTX2 U982 ( .A(n959), .B(n958), .Z(n960) );
  IVSVTX2 U983 ( .A(n1034), .Z(n1071) );
  IVSVTX6 U984 ( .A(n763), .Z(n673) );
  IVSVTX4 U985 ( .A(n990), .Z(n994) );
  OR2SVTX2 U986 ( .A(n310), .B(n970), .Z(n767) );
  IVSVTX2 U987 ( .A(n310), .Z(n606) );
  B_ND2SVTX2 U988 ( .A(N[0]), .B(n1003), .Z(n692) );
  IVSVTX2 U989 ( .A(n1003), .Z(n986) );
  CTIVSVTX2 U990 ( .A(n1280), .Z(n413) );
  ND2SVTX6 U991 ( .A(n549), .B(n548), .Z(n868) );
  CTIVSVTX2 U992 ( .A(n981), .Z(n412) );
  IVSVTX6 U993 ( .A(N[8]), .Z(n912) );
  AO7SVTX6 U994 ( .A(n1645), .B(n1644), .C(n1643), .Z(n1734) );
  B_ND2SVTX2 U995 ( .A(n1811), .B(n789), .Z(n1814) );
  OR2SVTX2 U996 ( .A(n1810), .B(n1809), .Z(n789) );
  IVSVTX2 U997 ( .A(n1721), .Z(n352) );
  IVSVTX4 U998 ( .A(n1641), .Z(n460) );
  IVSVTX4 U999 ( .A(n398), .Z(n1681) );
  IVSVTX2 U1000 ( .A(n1635), .Z(n434) );
  AO7ABSVTX6 U1001 ( .A(n1586), .B(n1585), .C(n339), .Z(n1635) );
  F_ENSVTX2 U1002 ( .A(n795), .B(n1616), .Z(n401) );
  ENSVTX4 U1003 ( .A(n1758), .B(n363), .Z(O[15]) );
  AO7SVTX2 U1004 ( .A(n1756), .B(n1759), .C(n1757), .Z(n363) );
  IVSVTX2 U1005 ( .A(n533), .Z(n532) );
  NR2SVTX2 U1006 ( .A(n1659), .B(n1658), .Z(n533) );
  AN2SVTX2 U1007 ( .A(n1612), .B(n1611), .Z(n795) );
  IVSVTX2 U1008 ( .A(n1660), .Z(n1662) );
  FAS1SVTX2 U1009 ( .A(n1629), .B(n616), .CI(n1428), .CO(n1651), .Z(n1637) );
  FAS1SVTX2 U1010 ( .A(n1603), .B(n1602), .CI(n1601), .CO(n1675), .Z(n1660) );
  IVSVTX4 U1011 ( .A(n694), .Z(n288) );
  B_ND2SVTX2 U1012 ( .A(n1438), .B(n1761), .Z(n1763) );
  IVSVTX4 U1013 ( .A(n1507), .Z(n1508) );
  AO7SVTX4 U1014 ( .A(n1229), .B(n1782), .C(n1780), .Z(n758) );
  B_ND2SVTX2 U1015 ( .A(n1773), .B(n1772), .Z(n1777) );
  ND3SVTX4 U1016 ( .A(n526), .B(n1556), .C(n1557), .Z(n525) );
  IVSVTX6 U1017 ( .A(n569), .Z(n1439) );
  NR2ASVTX6 U1018 ( .A(n1483), .B(n1482), .Z(n1490) );
  B_ND2SVTX1 U1019 ( .A(n1791), .B(n1790), .Z(n1795) );
  B_ND2SVTX2 U1020 ( .A(n1431), .B(n1430), .Z(n695) );
  ND2ASVTX6 U1021 ( .A(n1133), .B(n1227), .Z(n1780) );
  IVSVTX4 U1022 ( .A(n1803), .Z(n700) );
  ND2ASVTX6 U1023 ( .A(n348), .B(n1707), .Z(n349) );
  ND2SVTX4 U1024 ( .A(n365), .B(n364), .Z(n571) );
  IVSVTX4 U1025 ( .A(n1800), .Z(n290) );
  ND2SVTX4 U1026 ( .A(n341), .B(n342), .Z(n343) );
  NR2SVTX6 U1027 ( .A(n1458), .B(n427), .Z(n342) );
  ND3SVTX6 U1028 ( .A(n1195), .B(n1194), .C(n1196), .Z(n442) );
  ND3SVTX4 U1029 ( .A(n1540), .B(n1200), .C(n1191), .Z(n1192) );
  AO2SVTX6 U1030 ( .A(n1119), .B(n1235), .C(n1212), .D(n1402), .Z(n1173) );
  IVSVTX2 U1031 ( .A(n776), .Z(n644) );
  F_ENSVTX2 U1032 ( .A(n1182), .B(n1215), .Z(n747) );
  NR2SVTX4 U1033 ( .A(n1142), .B(n1808), .Z(n1225) );
  CTIVSVTX4 U1034 ( .A(n635), .Z(n610) );
  ND3SVTX4 U1035 ( .A(n1209), .B(n360), .C(n1200), .Z(n361) );
  NR2SVTX4 U1036 ( .A(n1538), .B(n1537), .Z(n1543) );
  IVSVTX8 U1037 ( .A(n660), .Z(n346) );
  IVSVTX4 U1038 ( .A(n1677), .Z(n1546) );
  AO7SVTX4 U1039 ( .A(n1536), .B(n556), .C(n1535), .Z(n1537) );
  ND4ABSVTX6 U1040 ( .A(n1392), .B(n1375), .C(n1373), .D(n1374), .Z(n1379) );
  IVSVTX8 U1041 ( .A(n1585), .Z(n295) );
  IVSVTX4 U1042 ( .A(n1376), .Z(n297) );
  ND3SVTX6 U1043 ( .A(n1530), .B(n1311), .C(n1310), .Z(n1677) );
  ND2SVTX4 U1044 ( .A(n567), .B(n509), .Z(n1322) );
  ND2ASVTX4 U1045 ( .A(O[27]), .B(n665), .Z(n1242) );
  ND2ASVTX6 U1046 ( .A(n597), .B(n1408), .Z(n1449) );
  IVSVTX2 U1047 ( .A(n1342), .Z(n1345) );
  IVSVTX2 U1048 ( .A(n1203), .Z(n301) );
  ND2SVTX4 U1049 ( .A(n1127), .B(n1128), .Z(n665) );
  ND2SVTX4 U1050 ( .A(n386), .B(n404), .Z(n1011) );
  AO7SVTX6 U1051 ( .A(n1309), .B(n1308), .C(n1307), .Z(n1532) );
  NR2ASVTX4 U1052 ( .A(n463), .B(n500), .Z(n1168) );
  AO7SVTX4 U1053 ( .A(n1035), .B(n1106), .C(n480), .Z(n1054) );
  AO7SVTX6 U1054 ( .A(n422), .B(n421), .C(n419), .Z(n489) );
  NR2SVTX4 U1055 ( .A(n1074), .B(n897), .Z(n1080) );
  IVSVTX4 U1056 ( .A(n953), .Z(n478) );
  ND3ASVTX6 U1057 ( .A(n418), .B(n1048), .C(n420), .Z(n419) );
  IVSVTX6 U1058 ( .A(n950), .Z(n664) );
  B_ND2SVTX2 U1059 ( .A(n1314), .B(n1276), .Z(n770) );
  IVSVTX4 U1060 ( .A(n653), .Z(n1013) );
  NR2SVTX4 U1061 ( .A(n1009), .B(n335), .Z(n749) );
  IVSVTX10 U1062 ( .A(n592), .Z(n1339) );
  ND3SVTX6 U1063 ( .A(n767), .B(n973), .C(n264), .Z(n1352) );
  NR2SVTX4 U1064 ( .A(n1180), .B(n1070), .Z(n336) );
  ND2SVTX6 U1065 ( .A(O[29]), .B(n1033), .Z(n397) );
  AO6SVTX4 U1066 ( .A(n1061), .B(n873), .C(n1000), .Z(n376) );
  ND3SVTX4 U1067 ( .A(n329), .B(n327), .C(n935), .Z(n1303) );
  IVSVTX12 U1068 ( .A(n1340), .Z(n306) );
  ND2SVTX6 U1069 ( .A(n852), .B(n949), .Z(n671) );
  IVSVTX6 U1070 ( .A(n957), .Z(n1070) );
  IVSVTX10 U1071 ( .A(n1010), .Z(n852) );
  NR2SVTX2 U1072 ( .A(n892), .B(n1071), .Z(n390) );
  IVSVTX2 U1073 ( .A(n1328), .Z(n1297) );
  NR3ABSVTX6 U1074 ( .A(n925), .B(n319), .C(n697), .Z(n952) );
  IVSVTX2 U1075 ( .A(n659), .Z(n658) );
  IVSVTX4 U1076 ( .A(n982), .Z(n450) );
  NR2SVTX6 U1077 ( .A(n993), .B(n994), .Z(n995) );
  IVSVTX2 U1078 ( .A(n799), .Z(n468) );
  ND2SVTX6 U1079 ( .A(n1061), .B(n1062), .Z(n1033) );
  IVSVTX2 U1080 ( .A(n798), .Z(n1287) );
  IVSVTX8 U1081 ( .A(n673), .Z(n674) );
  IVSVTX2 U1082 ( .A(n886), .Z(n887) );
  IVSVTX1 U1083 ( .A(n867), .Z(n516) );
  B_ND2SVTX2 U1084 ( .A(n1020), .B(n484), .Z(n1021) );
  ND2SVTX6 U1085 ( .A(n880), .B(n879), .Z(n520) );
  AO7ABSVTX2 U1086 ( .A(n812), .B(n1020), .C(n811), .Z(n816) );
  IVSVTX2 U1087 ( .A(n1006), .Z(n311) );
  ND2SVTX6 U1088 ( .A(n667), .B(n808), .Z(n809) );
  IVSVTX6 U1089 ( .A(N[2]), .Z(n1031) );
  CTIVSVTX6 U1090 ( .A(n313), .Z(n1112) );
  NR2SVTX6 U1091 ( .A(n1114), .B(n314), .Z(n1320) );
  ND2SVTX4 U1092 ( .A(n315), .B(n1112), .Z(n314) );
  ND2SVTX4 U1093 ( .A(n1108), .B(n1029), .Z(n313) );
  IVSVTX6 U1094 ( .A(N[24]), .Z(n650) );
  IVSVTX8 U1095 ( .A(n1606), .Z(n1722) );
  ND2SVTX4 U1096 ( .A(n1406), .B(n1455), .Z(n668) );
  ND3ABSVTX4 U1097 ( .A(n1060), .B(n892), .C(n974), .Z(n1455) );
  AO6SVTX6 U1098 ( .A(n551), .B(n1626), .C(n1624), .Z(n1627) );
  IVSVTX8 U1099 ( .A(N[26]), .Z(n863) );
  IVSVTX6 U1100 ( .A(n587), .Z(n958) );
  ND3SVTX8 U1101 ( .A(n1368), .B(n318), .C(n1369), .Z(n1398) );
  ND2SVTX4 U1102 ( .A(n1367), .B(n1366), .Z(n318) );
  AO7SVTX8 U1103 ( .A(n1177), .B(n701), .C(n1313), .Z(n1007) );
  IVSVTX2 U1104 ( .A(n1632), .Z(n1717) );
  IVSVTX12 U1105 ( .A(n306), .Z(n497) );
  ND2SVTX6 U1106 ( .A(n1681), .B(n1680), .Z(n1723) );
  ND2SVTX6 U1107 ( .A(n392), .B(n391), .Z(n378) );
  AO2SVTX8 U1108 ( .A(n974), .B(n1139), .C(n1366), .D(n395), .Z(n975) );
  AO3SVTX6 U1109 ( .A(n442), .B(n1197), .C(n488), .D(n690), .Z(n1206) );
  NR4ABSVTX8 U1110 ( .A(n928), .B(n650), .C(n838), .D(n837), .Z(n842) );
  ND3SVTX8 U1111 ( .A(n924), .B(n680), .C(n902), .Z(n838) );
  ND2SVTX4 U1112 ( .A(n1520), .B(n1522), .Z(n324) );
  AO7SVTX2 U1113 ( .A(n1341), .B(n565), .C(n1403), .Z(n1342) );
  NR3ABSVTX8 U1114 ( .A(n1201), .B(n1186), .C(n699), .Z(n1800) );
  ND2ASVTX8 U1115 ( .A(n1574), .B(n1604), .Z(n443) );
  NR2SVTX4 U1116 ( .A(n285), .B(n1396), .Z(n638) );
  ND2SVTX4 U1117 ( .A(n1596), .B(n326), .Z(n1643) );
  NR2SVTX6 U1118 ( .A(n1596), .B(n326), .Z(n1645) );
  ENSVTX8 U1119 ( .A(n436), .B(n435), .Z(n326) );
  IVSVTX10 U1120 ( .A(n1072), .Z(n722) );
  ND2SVTX8 U1121 ( .A(n943), .B(n1017), .Z(n1072) );
  AO6SVTX4 U1122 ( .A(n724), .B(n1278), .C(n936), .Z(n329) );
  IVSVTX10 U1123 ( .A(n330), .Z(n849) );
  ND2SVTX8 U1124 ( .A(n331), .B(n1030), .Z(n330) );
  NR2SVTX4 U1125 ( .A(n330), .B(n869), .Z(n805) );
  NR2SVTX6 U1126 ( .A(N[23]), .B(N[22]), .Z(n331) );
  IVSVTX4 U1127 ( .A(n335), .Z(n1177) );
  AO7SVTX6 U1128 ( .A(n646), .B(n334), .C(n333), .Z(n335) );
  ND2SVTX4 U1129 ( .A(n1031), .B(n646), .Z(n333) );
  IVSVTX4 U1130 ( .A(n356), .Z(n957) );
  NR2SVTX2 U1131 ( .A(n336), .B(n749), .Z(n404) );
  IVSVTX4 U1132 ( .A(n337), .Z(n1752) );
  AO6ASVTX1 U1133 ( .A(n1699), .B(n1485), .C(n337), .Z(n1759) );
  AO7ABSVTX8 U1134 ( .A(n1460), .B(n299), .C(n343), .Z(n1481) );
  ND2ASVTX8 U1135 ( .A(n345), .B(n344), .Z(n1160) );
  ND2SVTX4 U1136 ( .A(n741), .B(n920), .Z(n345) );
  ND2SVTX4 U1137 ( .A(n1211), .B(n346), .Z(n1194) );
  ND2SVTX4 U1138 ( .A(n301), .B(n346), .Z(n663) );
  ND2SVTX4 U1139 ( .A(n265), .B(n346), .Z(n476) );
  ND2SVTX4 U1140 ( .A(n346), .B(n747), .Z(n1185) );
  AO2SVTX2 U1141 ( .A(n1183), .B(n346), .C(n1163), .D(n1161), .Z(n1164) );
  AO7SVTX8 U1142 ( .A(n349), .B(n1701), .C(n1703), .Z(n1774) );
  ND2SVTX8 U1143 ( .A(n924), .B(n350), .Z(n870) );
  NR2SVTX8 U1144 ( .A(N[19]), .B(N[24]), .Z(n350) );
  AO7ABSVTX8 U1145 ( .A(n1636), .B(n1635), .C(n351), .Z(n1641) );
  AO7ABSVTX6 U1146 ( .A(n434), .B(n433), .C(n435), .Z(n351) );
  AO7SVTX6 U1147 ( .A(n1617), .B(n1716), .C(n293), .Z(n435) );
  B_ND2SVTX2 U1148 ( .A(n282), .B(n765), .Z(n353) );
  ND2SVTX2 U1149 ( .A(n1717), .B(n1716), .Z(n354) );
  ND2ASVTX6 U1150 ( .A(n1478), .B(n1145), .Z(n1224) );
  ND2SVTX8 U1151 ( .A(n356), .B(n852), .Z(n355) );
  AO6ABSVTX8 U1152 ( .A(n752), .B(n824), .C(n1075), .Z(n356) );
  ND2SVTX6 U1153 ( .A(n358), .B(n954), .Z(n575) );
  ND3SVTX8 U1154 ( .A(n762), .B(n1525), .C(n938), .Z(n358) );
  ND2SVTX4 U1155 ( .A(n358), .B(n788), .Z(n1588) );
  ND4ABSVTX8 U1156 ( .A(n664), .B(n953), .C(n358), .D(n1095), .Z(n939) );
  ND2SVTX6 U1157 ( .A(n1173), .B(n1172), .Z(n359) );
  ND2SVTX6 U1158 ( .A(n283), .B(n359), .Z(n1703) );
  NR2ASVTX8 U1159 ( .A(n300), .B(n359), .Z(n1701) );
  AO3SVTX6 U1160 ( .A(n242), .B(n1209), .C(n362), .D(n361), .Z(n1202) );
  IVSVTX4 U1161 ( .A(n643), .Z(n1200) );
  IVSVTX12 U1162 ( .A(n709), .Z(n1119) );
  NR3SVTX8 U1163 ( .A(n1170), .B(n1230), .C(n1256), .Z(n366) );
  IVSVTX4 U1164 ( .A(N[21]), .Z(n922) );
  AO7CSVTX6 U1165 ( .A(n1798), .B(n367), .C(n1444), .Z(n1770) );
  IVSVTX4 U1166 ( .A(n218), .Z(n1798) );
  ND2SVTX8 U1167 ( .A(n1018), .B(n368), .Z(n1022) );
  ND3ABSVTX8 U1168 ( .A(n861), .B(n368), .C(n860), .Z(n944) );
  ND3ABSVTX8 U1169 ( .A(n823), .B(n368), .C(n860), .Z(n990) );
  ND2ASVTX8 U1170 ( .A(n1072), .B(n737), .Z(n1073) );
  ND2ASVTX8 U1171 ( .A(n1665), .B(n1657), .Z(n461) );
  ND2SVTX8 U1172 ( .A(n461), .B(n1663), .Z(n1683) );
  NR2SVTX8 U1173 ( .A(n1560), .B(n1563), .Z(n1570) );
  NR2ASVTX8 U1174 ( .A(n294), .B(n1630), .Z(n1563) );
  NR2ASVTX8 U1175 ( .A(n1513), .B(n1607), .Z(n1560) );
  NR2SVTX8 U1176 ( .A(n1610), .B(n370), .Z(n1620) );
  NR2ASVTX8 U1177 ( .A(n1547), .B(n1599), .Z(n1610) );
  ND2SVTX6 U1178 ( .A(n1570), .B(n1569), .Z(n1591) );
  NR3SVTX8 U1179 ( .A(n1512), .B(n371), .C(n288), .Z(n1569) );
  ND3SVTX6 U1180 ( .A(n295), .B(n521), .C(n593), .Z(n373) );
  ND2SVTX8 U1181 ( .A(n372), .B(n445), .Z(n1606) );
  IVSVTX6 U1182 ( .A(n768), .Z(n372) );
  AO5ASVTX8 U1183 ( .B(n432), .A(n1660), .C(n444), .Z(n768) );
  AO17ASVTX8 U1184 ( .A(n295), .B(n1579), .C(n1506), .D(n373), .Z(n1511) );
  NR2SVTX4 U1185 ( .A(n375), .B(n374), .Z(n1086) );
  ND3SVTX6 U1186 ( .A(n1146), .B(n1149), .C(n1081), .Z(n374) );
  ND3ASVTX6 U1187 ( .A(n722), .B(n1139), .C(n256), .Z(n1146) );
  ND2ASVTX8 U1188 ( .A(n1361), .B(n1324), .Z(n1084) );
  ND2SVTX4 U1189 ( .A(n1124), .B(n377), .Z(n1085) );
  ND2ASVTX8 U1190 ( .A(n309), .B(n1036), .Z(n1139) );
  AN2SVTX6 U1191 ( .A(n1082), .B(n719), .Z(n773) );
  EO3SVTX8 U1192 ( .A(n281), .B(n393), .C(n378), .Z(n544) );
  ND2SVTX4 U1193 ( .A(n1582), .B(n384), .Z(n380) );
  IVSVTX4 U1194 ( .A(n1745), .Z(n381) );
  IVSVTX4 U1195 ( .A(n1642), .Z(n1644) );
  BFSVTX6 U1196 ( .A(n494), .Z(n385) );
  ND2SVTX8 U1197 ( .A(n911), .B(n656), .Z(n387) );
  ND2ASVTX8 U1198 ( .A(n986), .B(n387), .Z(n1009) );
  ND2SVTX6 U1199 ( .A(n296), .B(n388), .Z(n647) );
  IVSVTX4 U1200 ( .A(n393), .Z(n1638) );
  AO2SVTX6 U1201 ( .A(n1125), .B(n1124), .C(n1525), .D(n1126), .Z(n1127) );
  ND2SVTX4 U1202 ( .A(n1333), .B(n1332), .Z(n395) );
  ND2SVTX4 U1203 ( .A(n587), .B(n396), .Z(n1062) );
  ND2SVTX2 U1204 ( .A(n396), .B(n1292), .Z(n873) );
  ND3ASVTX6 U1205 ( .A(n852), .B(n397), .C(n1121), .Z(n480) );
  AO2SVTX2 U1206 ( .A(n1646), .B(n1631), .C(n1574), .D(n1632), .Z(n400) );
  NR2ASVTX8 U1207 ( .A(n1618), .B(n1640), .Z(n1732) );
  MUX21NSVTX4 U1208 ( .A(n311), .B(n276), .S(n1019), .Z(n701) );
  ND2SVTX4 U1209 ( .A(n1175), .B(n451), .Z(n1004) );
  ND2ASVTX8 U1210 ( .A(n402), .B(n895), .Z(n1175) );
  IVSVTX4 U1211 ( .A(n1166), .Z(n402) );
  IVSVTX12 U1212 ( .A(n948), .Z(n985) );
  NR2ASVTX2 U1213 ( .A(n720), .B(n587), .Z(n774) );
  ND2SVTX4 U1214 ( .A(n1185), .B(n1184), .Z(n699) );
  ND2SVTX4 U1215 ( .A(n1183), .B(n746), .Z(n1184) );
  ND2SVTX4 U1216 ( .A(n1567), .B(n1620), .Z(n1571) );
  IVSVTX8 U1217 ( .A(n437), .Z(n641) );
  NR2SVTX4 U1218 ( .A(n928), .B(n759), .Z(n821) );
  ND3SVTX8 U1219 ( .A(n961), .B(n960), .C(n522), .Z(n962) );
  IVSVTX2 U1220 ( .A(n312), .Z(n1003) );
  NR2SVTX6 U1221 ( .A(n870), .B(n869), .Z(n846) );
  AO7CSVTX8 U1222 ( .A(n1451), .B(n295), .C(n1478), .Z(n1416) );
  NR3SVTX6 U1223 ( .A(n1070), .B(n1446), .C(n1447), .Z(n1467) );
  IVSVTX0H U1224 ( .A(n1467), .Z(n1456) );
  CTBUFSVTX8 U1225 ( .A(n576), .Z(n471) );
  ND2SVTX4 U1226 ( .A(n308), .B(n950), .Z(n406) );
  IVSVTX4 U1227 ( .A(n1365), .Z(n408) );
  ND3SVTX4 U1228 ( .A(n360), .B(n1155), .C(n1200), .Z(n1193) );
  ND3SVTX8 U1229 ( .A(n1193), .B(n476), .C(n1192), .Z(n1210) );
  NR2SVTX4 U1230 ( .A(n1591), .B(n1571), .Z(n1572) );
  AO7ASVTX4 U1231 ( .A(n530), .B(n1623), .C(n1613), .Z(n1614) );
  BFSVTX1 U1232 ( .A(n1476), .Z(n411) );
  AO6SVTX8 U1233 ( .A(n1716), .B(n1717), .C(n541), .Z(n1633) );
  AO7CSVTX4 U1234 ( .A(n1621), .B(n1623), .C(n1622), .Z(n1624) );
  NR2SVTX6 U1235 ( .A(N[24]), .B(N[26]), .Z(n414) );
  NR3ABSVTX8 U1236 ( .A(n659), .B(n416), .C(n1447), .Z(n1405) );
  IVSVTX4 U1237 ( .A(n306), .Z(n416) );
  AO7SVTX8 U1238 ( .A(n1045), .B(n417), .C(n1016), .Z(n1105) );
  NR2SVTX8 U1239 ( .A(n1083), .B(n309), .Z(n1046) );
  ND2ASVTX6 U1240 ( .A(n888), .B(n1294), .Z(n1039) );
  IVSVTX4 U1241 ( .A(n422), .Z(n1049) );
  ND2SVTX4 U1242 ( .A(n722), .B(n1040), .Z(n1048) );
  ND2SVTX4 U1243 ( .A(n1051), .B(n1050), .Z(n421) );
  IVSVTX4 U1244 ( .A(n875), .Z(n1058) );
  ND2SVTX4 U1245 ( .A(n722), .B(n1123), .Z(n1051) );
  ND2ASVTX8 U1246 ( .A(n423), .B(n1019), .Z(n422) );
  AO6ASVTX8 U1247 ( .A(n425), .B(n774), .C(n450), .Z(n1023) );
  AN2SVTX4 U1248 ( .A(n312), .B(n1022), .Z(n425) );
  IVSVTX4 U1249 ( .A(n1037), .Z(n426) );
  ND2ASVTX8 U1250 ( .A(n515), .B(n1017), .Z(n1037) );
  IVSVTX4 U1251 ( .A(n1481), .Z(n1479) );
  IVSVTX4 U1252 ( .A(n1470), .Z(n427) );
  ND2SVTX4 U1253 ( .A(n772), .B(n428), .Z(n1460) );
  F_ENSVTX2 U1254 ( .A(n1519), .B(n1518), .Z(n431) );
  F_ENSVTX2 U1255 ( .A(n1636), .B(n1635), .Z(n436) );
  AO7ABSVTX8 U1256 ( .A(n1603), .B(n449), .C(n1382), .Z(n1384) );
  AO7SVTX6 U1257 ( .A(n1736), .B(n1732), .C(n438), .Z(n487) );
  ND2SVTX1 U1258 ( .A(n438), .B(n1733), .Z(n1738) );
  ND2SVTX8 U1259 ( .A(n803), .B(n439), .Z(n675) );
  NR2SVTX6 U1260 ( .A(N[17]), .B(N[16]), .Z(n439) );
  IVSVTX6 U1261 ( .A(N[27]), .Z(n803) );
  IVSVTX4 U1262 ( .A(n878), .Z(n440) );
  ND2SVTX6 U1263 ( .A(n944), .B(n440), .Z(n754) );
  NR2SVTX4 U1264 ( .A(N[20]), .B(N[22]), .Z(n832) );
  ND2SVTX4 U1265 ( .A(n1197), .B(n442), .Z(n1207) );
  IVSVTX4 U1266 ( .A(n1661), .Z(n444) );
  ND2SVTX8 U1267 ( .A(n689), .B(n1018), .Z(n448) );
  NR3ABSVTX8 U1268 ( .A(n826), .B(n849), .C(n448), .Z(n867) );
  IVSVTX4 U1269 ( .A(n1542), .Z(n449) );
  ND2SVTX8 U1270 ( .A(n1292), .B(n889), .Z(n1036) );
  BFSVTX8 U1271 ( .A(N[22]), .Z(n901) );
  ND2SVTX4 U1272 ( .A(n1003), .B(n1082), .Z(n452) );
  ND2SVTX8 U1273 ( .A(n962), .B(n576), .Z(n1249) );
  NR3ABSVTX8 U1274 ( .A(n1020), .B(n872), .C(n462), .Z(n979) );
  IVSVTX8 U1275 ( .A(n1356), .Z(n1365) );
  ND3ABSVTX6 U1276 ( .A(n872), .B(n276), .C(n752), .Z(n1015) );
  AO7SVTX8 U1277 ( .A(n289), .B(n1219), .C(n1218), .Z(n1435) );
  ND2SVTX6 U1278 ( .A(n1049), .B(n514), .Z(n1103) );
  ND3SVTX8 U1279 ( .A(n1542), .B(n1547), .C(n1555), .Z(n1382) );
  MUX21NSVTX6 U1280 ( .A(n1396), .B(n1534), .S(n500), .Z(n1318) );
  NR2SVTX4 U1281 ( .A(n1701), .B(n1174), .Z(n1775) );
  ENSVTX8 U1282 ( .A(n458), .B(n457), .Z(n1680) );
  F_ENSVTX2 U1283 ( .A(n1720), .B(n1719), .Z(n458) );
  ND3SVTX8 U1284 ( .A(n851), .B(n850), .C(n459), .Z(n983) );
  ND2ASVTX8 U1285 ( .A(n460), .B(n544), .Z(n1736) );
  IVSVTX12 U1286 ( .A(n1604), .Z(n1716) );
  IVSVTX6 U1287 ( .A(n948), .Z(n1106) );
  BFSVTX12 U1288 ( .A(n1017), .Z(n462) );
  AO17SVTX8 U1289 ( .A(n1504), .B(n1503), .C(n1502), .D(n786), .Z(n1625) );
  ND3SVTX8 U1290 ( .A(n1436), .B(n1693), .C(n1435), .Z(n1504) );
  ND2SVTX4 U1291 ( .A(n1364), .B(n1522), .Z(n1369) );
  AO6SVTX8 U1292 ( .A(n1625), .B(n1577), .C(n465), .Z(n1578) );
  AO7SVTX8 U1293 ( .A(n1576), .B(n1623), .C(n735), .Z(n465) );
  ND3ABSVTX8 U1294 ( .A(n634), .B(n1513), .C(n559), .Z(n557) );
  ND4SVTX8 U1295 ( .A(n1002), .B(n1154), .C(n561), .D(n648), .Z(n736) );
  AO2SVTX4 U1296 ( .A(n306), .B(n997), .C(n1340), .D(n996), .Z(n684) );
  ND3SVTX8 U1297 ( .A(n964), .B(n912), .C(n810), .Z(n672) );
  MUX21NSVTX8 U1298 ( .A(n997), .B(n1023), .S(n743), .Z(n1100) );
  IVSVTX12 U1299 ( .A(n1082), .Z(n1124) );
  ND2SVTX8 U1300 ( .A(n1649), .B(n275), .Z(n545) );
  NR3ABSVTX4 U1301 ( .A(N[21]), .B(n941), .C(n822), .Z(n819) );
  ND2SVTX8 U1302 ( .A(n944), .B(n535), .Z(n910) );
  IVSVTX6 U1303 ( .A(n489), .Z(n1052) );
  ND3SVTX8 U1304 ( .A(n466), .B(n976), .C(n975), .Z(n1343) );
  ND2SVTX4 U1305 ( .A(n1352), .B(n1324), .Z(n466) );
  NR2ASVTX2 U1306 ( .A(N[1]), .B(n752), .Z(n971) );
  ND2ASVTX8 U1307 ( .A(n712), .B(n536), .Z(n521) );
  NR2SVTX4 U1308 ( .A(n952), .B(n565), .Z(n496) );
  ND2SVTX4 U1309 ( .A(n469), .B(n468), .Z(n653) );
  BFSVTX1 U1310 ( .A(n1405), .Z(n472) );
  IVSVTX4 U1311 ( .A(n752), .Z(n473) );
  NR2SVTX4 U1312 ( .A(n473), .B(n874), .Z(n875) );
  IVSVTX4 U1313 ( .A(n474), .Z(n788) );
  ND2SVTX4 U1314 ( .A(n478), .B(n1095), .Z(n474) );
  ND2SVTX8 U1315 ( .A(n782), .B(n1731), .Z(n1741) );
  BFSVTX2 U1316 ( .A(n1188), .Z(n475) );
  NR3SVTX6 U1317 ( .A(n1255), .B(n1256), .C(n1264), .Z(n1153) );
  NR4ABCSVTX6 U1318 ( .A(n1338), .B(n625), .C(n1407), .D(n1337), .Z(n1346) );
  ND2SVTX6 U1319 ( .A(n1781), .B(n1711), .Z(n1238) );
  IVSVTX6 U1320 ( .A(N[25]), .Z(n928) );
  NR2SVTX6 U1321 ( .A(n267), .B(n590), .Z(n1241) );
  ND3SVTX8 U1322 ( .A(n651), .B(n315), .C(n1112), .Z(n1056) );
  IVSVTX8 U1323 ( .A(n1285), .Z(n932) );
  IVSVTX4 U1324 ( .A(n845), .Z(n807) );
  NR2SVTX4 U1325 ( .A(n1398), .B(n1412), .Z(n1374) );
  ND2SVTX4 U1326 ( .A(n1363), .B(n1362), .Z(n1412) );
  ND3ASVTX6 U1327 ( .A(n479), .B(n1221), .C(n572), .Z(n485) );
  IVSVTX4 U1328 ( .A(n1262), .Z(n1135) );
  ND3ABSVTX8 U1329 ( .A(n1416), .B(n482), .C(n481), .Z(n1421) );
  IVSVTX8 U1330 ( .A(n546), .Z(n559) );
  ND2SVTX4 U1331 ( .A(n601), .B(n305), .Z(n1147) );
  ND4SVTX6 U1332 ( .A(N[7]), .B(n861), .C(n928), .D(n677), .Z(n833) );
  ENSVTX8 U1333 ( .A(n1470), .B(n1264), .Z(n1145) );
  IVSVTX4 U1334 ( .A(n924), .Z(n760) );
  ND4SVTX6 U1335 ( .A(n829), .B(n761), .C(n723), .D(n849), .Z(n830) );
  AO3NSVTX8 U1336 ( .A(n1752), .B(n1501), .C(n1500), .D(n1750), .Z(n786) );
  IVSVTX2 U1337 ( .A(n1464), .Z(n1465) );
  ND2ASVTX8 U1338 ( .A(n601), .B(n1343), .Z(n1067) );
  ND2SVTX4 U1339 ( .A(n949), .B(n852), .Z(n921) );
  ND2ASVTX8 U1340 ( .A(n1057), .B(n284), .Z(n1170) );
  ND2SVTX4 U1341 ( .A(n491), .B(n1246), .Z(n1078) );
  ND2SVTX4 U1342 ( .A(n1077), .B(n492), .Z(n491) );
  AO7SVTX6 U1343 ( .A(n1132), .B(n266), .C(n693), .Z(n1262) );
  IVSVTX8 U1344 ( .A(n983), .Z(n656) );
  F_ENSVTX2 U1345 ( .A(n1182), .B(n1215), .Z(n1191) );
  IVSVTX4 U1346 ( .A(n493), .Z(n1182) );
  ND4ABSVTX8 U1347 ( .A(n385), .B(n1181), .C(n265), .D(n511), .Z(n493) );
  ND2SVTX4 U1348 ( .A(n1801), .B(n495), .Z(n1705) );
  ND2SVTX4 U1349 ( .A(n700), .B(n290), .Z(n495) );
  IVSVTX6 U1350 ( .A(n618), .Z(n541) );
  AO2SVTX6 U1351 ( .A(n585), .B(n636), .C(n1398), .D(O[27]), .Z(n626) );
  NR2SVTX4 U1352 ( .A(n953), .B(n496), .Z(n954) );
  ND2SVTX4 U1353 ( .A(n307), .B(n1523), .Z(n920) );
  ND2SVTX4 U1354 ( .A(n1025), .B(n1024), .Z(n498) );
  IVSVTX8 U1355 ( .A(n1340), .Z(n1043) );
  IVSVTX4 U1356 ( .A(n1525), .Z(O[28]) );
  IVSVTX8 U1357 ( .A(n763), .Z(n1292) );
  BFSVTX6 U1358 ( .A(n1140), .Z(n500) );
  ND3SVTX8 U1359 ( .A(n964), .B(n912), .C(n810), .Z(n856) );
  EOSVTX8 U1360 ( .A(n619), .B(n1401), .Z(n540) );
  ND2ASVTX8 U1361 ( .A(n1513), .B(n1607), .Z(n1562) );
  ND2SVTX4 U1362 ( .A(n1749), .B(n598), .Z(n1500) );
  ND4ABSVTX8 U1363 ( .A(n1499), .B(n600), .C(n599), .D(n1497), .Z(n1749) );
  IVSVTX12 U1364 ( .A(n584), .Z(n1340) );
  ENSVTX8 U1365 ( .A(n1652), .B(n537), .Z(n536) );
  ND3SVTX6 U1366 ( .A(n1144), .B(n1221), .C(n572), .Z(n1711) );
  ND2SVTX6 U1367 ( .A(n1652), .B(n1630), .Z(n1561) );
  ND2SVTX4 U1368 ( .A(n1367), .B(n1365), .Z(n1330) );
  IVSVTX4 U1369 ( .A(n1452), .Z(n1458) );
  B_ND2SVTX2 U1370 ( .A(n296), .B(n1119), .Z(n776) );
  NR3ABSVTX2 U1371 ( .A(N[3]), .B(n484), .C(n853), .Z(n799) );
  ND2ASVTX8 U1372 ( .A(n985), .B(n583), .Z(n1111) );
  IVSVTX4 U1373 ( .A(n1190), .Z(n1094) );
  ND2SVTX4 U1374 ( .A(n1305), .B(n1306), .Z(n503) );
  BFSVTX4 U1375 ( .A(N[14]), .Z(n940) );
  AO7ABSVTX4 U1376 ( .A(n1023), .B(n1340), .C(n652), .Z(n1108) );
  ND3ABSVTX8 U1377 ( .A(n909), .B(n867), .C(n656), .Z(n1010) );
  IVSVTX12 U1378 ( .A(n646), .Z(n1019) );
  IVSVTX8 U1379 ( .A(n563), .Z(n1092) );
  ND3SVTX6 U1380 ( .A(n726), .B(n505), .C(n858), .Z(n943) );
  ND2ASVTX8 U1381 ( .A(n757), .B(n1421), .Z(n604) );
  ND2SVTX4 U1382 ( .A(n1209), .B(n1208), .Z(n1801) );
  AO6SVTX8 U1383 ( .A(n1305), .B(n1306), .C(n1073), .Z(n953) );
  ND3SVTX6 U1384 ( .A(n507), .B(n1321), .C(n508), .Z(n1323) );
  IVSVTX4 U1385 ( .A(n1322), .Z(n507) );
  ND2ASVTX8 U1386 ( .A(n984), .B(n894), .Z(n646) );
  IVSVTX4 U1387 ( .A(n734), .Z(n511) );
  NR2SVTX4 U1388 ( .A(n1255), .B(n1256), .Z(n512) );
  ND2ASVTX8 U1389 ( .A(N[26]), .B(n1314), .Z(n837) );
  AO7ABSVTX8 U1390 ( .A(n1068), .B(n703), .C(n1067), .Z(n563) );
  ND2ASVTX8 U1391 ( .A(n818), .B(n1022), .Z(n853) );
  IVSVTX4 U1392 ( .A(n932), .Z(n724) );
  ND2ASVTX8 U1393 ( .A(n296), .B(n513), .Z(n1437) );
  OR2SVTX8 U1394 ( .A(n932), .B(n763), .Z(n1291) );
  ND2ASVTX8 U1395 ( .A(n514), .B(n579), .Z(n580) );
  ND3ABSVTX4 U1396 ( .A(n1720), .B(n717), .C(n1554), .Z(n1544) );
  ND3SVTX4 U1397 ( .A(n936), .B(n902), .C(n862), .Z(n839) );
  ND2SVTX4 U1398 ( .A(n1352), .B(n1522), .Z(n1407) );
  NR3SVTX6 U1399 ( .A(n678), .B(n1466), .C(n1255), .Z(n1093) );
  AO2SVTX6 U1400 ( .A(n1521), .B(n1365), .C(n1366), .D(n1364), .Z(n1298) );
  ND2SVTX4 U1401 ( .A(n742), .B(n1437), .Z(n1443) );
  ND2SVTX8 U1402 ( .A(n519), .B(n518), .Z(n1607) );
  AO2ABSVTX6 U1403 ( .C(n526), .D(n617), .A(n1808), .B(n1566), .Z(n519) );
  B_IVSVTX1 U1404 ( .A(n520), .Z(n817) );
  ND2SVTX4 U1405 ( .A(n593), .B(n521), .Z(n1579) );
  EO3SVTX8 U1406 ( .A(n1662), .B(n443), .C(n1661), .Z(n1666) );
  ND2ASVTX8 U1407 ( .A(n527), .B(n525), .Z(n1599) );
  IVSVTX4 U1408 ( .A(n753), .Z(n526) );
  AO17SVTX4 U1409 ( .A(n528), .B(n1558), .C(n745), .D(n1559), .Z(n527) );
  IVSVTX4 U1410 ( .A(n529), .Z(n528) );
  ND2SVTX4 U1411 ( .A(n1555), .B(n1542), .Z(n529) );
  ND4SVTX8 U1412 ( .A(n1566), .B(n1552), .C(n1551), .D(n1550), .Z(n530) );
  ND2SVTX6 U1413 ( .A(n1544), .B(n1545), .Z(n1551) );
  ND2SVTX8 U1414 ( .A(n1664), .B(n1665), .Z(n1739) );
  ENSVTX8 U1415 ( .A(n1653), .B(n545), .Z(n1665) );
  NR2ASVTX6 U1416 ( .A(n1667), .B(n1666), .Z(n531) );
  ND2ASVTX8 U1417 ( .A(n866), .B(n865), .Z(n878) );
  NR2SVTX8 U1418 ( .A(n867), .B(n878), .Z(n535) );
  NR3SVTX8 U1419 ( .A(n539), .B(n1428), .C(n538), .Z(n537) );
  ND3SVTX4 U1420 ( .A(n1418), .B(n1419), .C(n633), .Z(n538) );
  ND2ASVTX8 U1421 ( .A(n303), .B(n1399), .Z(n1428) );
  IVSVTX4 U1422 ( .A(n739), .Z(n539) );
  ND2SVTX4 U1423 ( .A(n1315), .B(n576), .Z(n542) );
  BFSVTX6 U1424 ( .A(n1574), .Z(n543) );
  ND2SVTX6 U1425 ( .A(n1728), .B(n286), .Z(n1730) );
  ND3SVTX8 U1426 ( .A(n1419), .B(n1418), .C(n739), .Z(n546) );
  NR2SVTX4 U1427 ( .A(n1585), .B(n546), .Z(n555) );
  AO7SVTX6 U1428 ( .A(n292), .B(n546), .C(n1513), .Z(n558) );
  ND2SVTX4 U1429 ( .A(n710), .B(n775), .Z(n1137) );
  ENSVTX0H U1430 ( .A(n551), .B(n1779), .Z(O[16]) );
  NR2SVTX6 U1431 ( .A(N[26]), .B(N[24]), .Z(n548) );
  ND2SVTX8 U1432 ( .A(n550), .B(n862), .Z(n818) );
  NR2SVTX8 U1433 ( .A(N[29]), .B(N[28]), .Z(n862) );
  NR2SVTX6 U1434 ( .A(N[31]), .B(N[30]), .Z(n550) );
  AO17SVTX8 U1435 ( .A(n1504), .B(n1503), .C(n1502), .D(n786), .Z(n551) );
  ND2SVTX6 U1436 ( .A(n552), .B(n553), .Z(n1495) );
  AO6SVTX8 U1437 ( .A(n654), .B(n1483), .C(n1462), .Z(n553) );
  IVSVTX4 U1438 ( .A(n1757), .Z(n598) );
  ND2SVTX8 U1439 ( .A(n1496), .B(n1495), .Z(n1757) );
  ND3ASVTX4 U1440 ( .A(n600), .B(n599), .C(n1497), .Z(n1498) );
  ND2SVTX8 U1441 ( .A(n560), .B(n554), .Z(n1497) );
  IVSVTX6 U1442 ( .A(n1420), .Z(n603) );
  ND2SVTX8 U1443 ( .A(n560), .B(n649), .Z(n1420) );
  ND2SVTX8 U1444 ( .A(n557), .B(n558), .Z(n649) );
  ND2SVTX6 U1445 ( .A(n987), .B(n1187), .Z(n561) );
  NR2SVTX4 U1446 ( .A(n1465), .B(n563), .Z(n1469) );
  ND2SVTX4 U1447 ( .A(n564), .B(n1092), .Z(n784) );
  IVSVTX4 U1448 ( .A(n1466), .Z(n564) );
  ND2ASVTX8 U1449 ( .A(n722), .B(n671), .Z(n681) );
  BFSVTX12 U1450 ( .A(n681), .Z(n565) );
  NR2ASVTX6 U1451 ( .A(n282), .B(n1479), .Z(n1461) );
  IVSVTX4 U1452 ( .A(n1057), .Z(n567) );
  ND2ASVTX8 U1453 ( .A(n685), .B(n568), .Z(n1057) );
  ND2SVTX4 U1454 ( .A(n1106), .B(n1156), .Z(n568) );
  ND2SVTX2 U1455 ( .A(n569), .B(n742), .Z(n1272) );
  ND2ASVTX8 U1456 ( .A(n1099), .B(n688), .Z(n569) );
  ND2SVTX4 U1457 ( .A(n962), .B(n1365), .Z(n968) );
  IVSVTX4 U1458 ( .A(n571), .Z(n1214) );
  ND2SVTX4 U1459 ( .A(n1216), .B(n571), .Z(n1772) );
  ND2SVTX4 U1460 ( .A(n1136), .B(n291), .Z(n572) );
  ND3SVTX8 U1461 ( .A(n574), .B(n1224), .C(n1226), .Z(n1227) );
  ND2SVTX8 U1462 ( .A(n1483), .B(n573), .Z(n1226) );
  ND2SVTX4 U1463 ( .A(n576), .B(n926), .Z(n1095) );
  NR2SVTX2 U1464 ( .A(n915), .B(n763), .Z(n577) );
  ND2SVTX4 U1465 ( .A(n1402), .B(n578), .Z(n645) );
  ENSVTX8 U1466 ( .A(n1258), .B(n1243), .Z(n578) );
  IVSVTX4 U1467 ( .A(n241), .Z(n581) );
  ND2SVTX8 U1468 ( .A(n995), .B(n656), .Z(n584) );
  ND3SVTX8 U1469 ( .A(n1353), .B(n1354), .C(n1355), .Z(n585) );
  AO2SVTX6 U1470 ( .A(n1414), .B(n556), .C(n1413), .D(n585), .Z(n1415) );
  IVSVTX12 U1471 ( .A(n586), .Z(n777) );
  IVSVTX12 U1472 ( .A(n872), .Z(n587) );
  ND2ASVTX8 U1473 ( .A(n872), .B(n885), .Z(n586) );
  ND2SVTX8 U1474 ( .A(n291), .B(n573), .Z(n588) );
  ND2SVTX6 U1475 ( .A(n1791), .B(n1237), .Z(n1712) );
  ND2ASVTX8 U1476 ( .A(n284), .B(n589), .Z(n1792) );
  ND3ASVTX8 U1477 ( .A(n792), .B(n687), .C(n686), .Z(n589) );
  ND2SVTX6 U1478 ( .A(n1241), .B(n1242), .Z(n1264) );
  ND2SVTX4 U1479 ( .A(n1141), .B(n666), .Z(n590) );
  ND3ABSVTX6 U1480 ( .A(n515), .B(n276), .C(n1017), .Z(n988) );
  AO6CSVTX8 U1481 ( .A(n649), .B(n291), .C(n1423), .Z(n593) );
  AO6ASVTX8 U1482 ( .A(n285), .B(n1449), .C(n594), .Z(n1452) );
  IVSVTX4 U1483 ( .A(n595), .Z(n594) );
  ND2SVTX4 U1484 ( .A(n625), .B(n1448), .Z(n596) );
  ND2SVTX4 U1485 ( .A(n1406), .B(n1407), .Z(n597) );
  ND2SVTX4 U1486 ( .A(n500), .B(n625), .Z(n790) );
  NR2ASVTX6 U1487 ( .A(n556), .B(n1394), .Z(n1395) );
  ND2SVTX4 U1488 ( .A(n556), .B(n1388), .Z(n714) );
  ND2SVTX6 U1489 ( .A(n1419), .B(n1418), .Z(n615) );
  ND2SVTX6 U1490 ( .A(n611), .B(n609), .Z(n1427) );
  ND3SVTX8 U1491 ( .A(n635), .B(n614), .C(n612), .Z(n611) );
  NR2SVTX8 U1492 ( .A(n1650), .B(n613), .Z(n612) );
  ND2SVTX6 U1493 ( .A(n1399), .B(n739), .Z(n613) );
  AO7SVTX8 U1494 ( .A(n1395), .B(n638), .C(n1397), .Z(n1650) );
  IVSVTX4 U1495 ( .A(n1427), .Z(n617) );
  ND2SVTX6 U1496 ( .A(n1339), .B(n1140), .Z(n620) );
  IVSVTX4 U1497 ( .A(n257), .Z(n622) );
  ND2SVTX8 U1498 ( .A(n623), .B(n1285), .Z(n725) );
  AO17ASVTX6 U1499 ( .A(n720), .B(n778), .C(n884), .D(n883), .Z(n623) );
  ND2SVTX4 U1500 ( .A(n969), .B(n1366), .Z(n625) );
  NR2SVTX6 U1501 ( .A(n629), .B(n1424), .Z(n635) );
  ND2SVTX6 U1502 ( .A(n285), .B(n1414), .Z(n628) );
  ND3SVTX4 U1503 ( .A(n637), .B(n714), .C(n630), .Z(n629) );
  NR3SVTX4 U1504 ( .A(n632), .B(n303), .C(n631), .Z(n630) );
  ND3SVTX6 U1505 ( .A(n714), .B(n637), .C(n297), .Z(n1652) );
  ND2SVTX6 U1506 ( .A(n639), .B(n640), .Z(n688) );
  ND2SVTX4 U1507 ( .A(n642), .B(n1164), .Z(n1707) );
  AO7SVTX8 U1508 ( .A(n1647), .B(n1427), .C(n1426), .Z(n1507) );
  NR2SVTX8 U1509 ( .A(n1190), .B(n643), .Z(n956) );
  ND2SVTX6 U1510 ( .A(n766), .B(n1097), .Z(n643) );
  IVSVTX6 U1511 ( .A(n647), .Z(n702) );
  IVSVTX4 U1512 ( .A(n499), .Z(n1169) );
  ND2SVTX6 U1513 ( .A(n1106), .B(n1100), .Z(n648) );
  NR2SVTX6 U1514 ( .A(n1105), .B(n1100), .Z(n651) );
  ND2SVTX4 U1515 ( .A(n1340), .B(n653), .Z(n1016) );
  ND2SVTX8 U1516 ( .A(n655), .B(n863), .Z(n845) );
  ND2SVTX4 U1517 ( .A(n659), .B(n1335), .Z(n1445) );
  ND2SVTX4 U1518 ( .A(n1333), .B(n1332), .Z(n659) );
  ND2SVTX6 U1519 ( .A(n766), .B(n1097), .Z(n955) );
  ND2ASVTX8 U1520 ( .A(n1190), .B(n955), .Z(n660) );
  IVSVTX4 U1521 ( .A(n856), .Z(n879) );
  NR2SVTX6 U1522 ( .A(N[15]), .B(N[13]), .Z(n667) );
  NR2SVTX4 U1523 ( .A(n809), .B(n856), .Z(n723) );
  NR2SVTX4 U1524 ( .A(n668), .B(n1068), .Z(n1348) );
  ND2SVTX4 U1525 ( .A(n1250), .B(n1249), .Z(n1068) );
  NR2SVTX4 U1526 ( .A(n670), .B(n669), .Z(n1431) );
  AO6SVTX4 U1527 ( .A(n1513), .B(n1429), .C(n294), .Z(n670) );
  ND4ABSVTX8 U1528 ( .A(n672), .B(n836), .C(n880), .D(n835), .Z(n851) );
  ND2SVTX8 U1529 ( .A(n310), .B(n885), .Z(n763) );
  ND2ASVTX8 U1530 ( .A(n1142), .B(n676), .Z(n1764) );
  ND2SVTX4 U1531 ( .A(n1198), .B(n332), .Z(n1203) );
  NR2SVTX4 U1532 ( .A(N[17]), .B(N[30]), .Z(n677) );
  IVSVTX4 U1533 ( .A(N[18]), .Z(n861) );
  NR2SVTX4 U1534 ( .A(n678), .B(n1170), .Z(n1171) );
  NR2SVTX8 U1535 ( .A(n678), .B(n1255), .Z(n1470) );
  ND2ASVTX8 U1536 ( .A(n1647), .B(n1267), .Z(n1268) );
  ND2SVTX8 U1537 ( .A(n1094), .B(n955), .Z(n1478) );
  ND2SVTX4 U1538 ( .A(n985), .B(n684), .Z(n1154) );
  ND2SVTX4 U1539 ( .A(n1525), .B(n685), .Z(n1157) );
  IVSVTX4 U1540 ( .A(n1792), .Z(n1236) );
  CTIVSVTX6 U1541 ( .A(n688), .Z(n1098) );
  IVSVTX4 U1542 ( .A(n838), .Z(n689) );
  IVSVTX4 U1543 ( .A(n698), .Z(n1304) );
  NR2SVTX4 U1544 ( .A(n1279), .B(n1291), .Z(n698) );
  ND2ASVTX8 U1545 ( .A(n1211), .B(n1210), .Z(n1803) );
  ND3SVTX4 U1546 ( .A(n1123), .B(n1122), .C(n949), .Z(n1077) );
  AO7SVTX2 U1547 ( .A(n1515), .B(n1514), .C(n1562), .Z(n1516) );
  ENSVTX8 U1548 ( .A(n1230), .B(n1171), .Z(n1212) );
  ND2SVTX2 U1549 ( .A(n1130), .B(n285), .Z(n1131) );
  AO7SVTX2 U1550 ( .A(n1526), .B(n1525), .C(n1524), .Z(n1587) );
  AO6ABSVTX6 U1551 ( .A(O[29]), .B(n1290), .C(n918), .Z(n1526) );
  ND3SVTX4 U1552 ( .A(n279), .B(n1555), .C(n1554), .Z(n1556) );
  MUX21NSVTX6 U1553 ( .A(n1251), .B(n1152), .S(n703), .Z(n900) );
  AO7ABSVTX4 U1554 ( .A(n996), .B(n355), .C(n1001), .Z(n1002) );
  IVSVTX8 U1555 ( .A(n355), .Z(n1387) );
  IVSVTX4 U1556 ( .A(n704), .Z(n705) );
  IVSVTX6 U1557 ( .A(N[30]), .Z(n902) );
  NR3SVTX4 U1558 ( .A(n906), .B(n905), .C(n904), .Z(n741) );
  IVSVTX12 U1559 ( .A(n1110), .Z(n1256) );
  AO7ABSVTX8 U1560 ( .A(n748), .B(n1370), .C(n1372), .Z(n1411) );
  ND2SVTX4 U1561 ( .A(n500), .B(n1388), .Z(n706) );
  NR2ASVTX2 U1562 ( .A(n1736), .B(n732), .Z(n1742) );
  AO7SVTX4 U1563 ( .A(n1722), .B(n1684), .C(n1724), .Z(n1685) );
  AO4ABSVTX6 U1564 ( .C(n1325), .D(n887), .A(n933), .B(n1294), .Z(n1370) );
  ND2SVTX4 U1565 ( .A(n969), .B(n748), .Z(n1363) );
  IVSVTX12 U1566 ( .A(n1350), .Z(n1542) );
  ND2ASVTX4 U1567 ( .A(n1467), .B(n1464), .Z(n1493) );
  ND2SVTX2 U1568 ( .A(n1523), .B(n1365), .Z(n1524) );
  ND3SVTX4 U1569 ( .A(n1280), .B(n674), .C(n724), .Z(n1281) );
  ND2SVTX4 U1570 ( .A(n962), .B(n748), .Z(n1390) );
  ND2ASVTX8 U1571 ( .A(n794), .B(n1812), .Z(n1813) );
  ND3SVTX8 U1572 ( .A(n731), .B(n1734), .C(n1733), .Z(n1731) );
  AO2SVTX2 U1573 ( .A(n1365), .B(n1315), .C(n1313), .D(n1314), .Z(n1529) );
  ND2SVTX4 U1574 ( .A(n1302), .B(n1301), .Z(n1534) );
  AO6SVTX2 U1575 ( .A(n282), .B(n1473), .C(n781), .Z(n1474) );
  NR2ASVTX2 U1576 ( .A(n530), .B(n1591), .Z(n1615) );
  ND3SVTX4 U1577 ( .A(n1075), .B(n1076), .C(n1339), .Z(n1246) );
  ND2ASVTX8 U1578 ( .A(n716), .B(n1573), .Z(n1574) );
  AO7SVTX2 U1579 ( .A(n1571), .B(n1623), .C(n1568), .Z(n716) );
  IVSVTX8 U1580 ( .A(n901), .Z(n941) );
  IVSVTX2 U1581 ( .A(n1040), .Z(n719) );
  IVSVTX4 U1582 ( .A(n1083), .Z(n1040) );
  IVSVTX4 U1583 ( .A(n731), .Z(n732) );
  ND2SVTX4 U1584 ( .A(n1258), .B(n1119), .Z(n1259) );
  ENSVTX8 U1585 ( .A(n1476), .B(n1093), .Z(n1267) );
  ND2SVTX2 U1586 ( .A(n950), .B(n1534), .Z(n1311) );
  AO6SVTX4 U1587 ( .A(n817), .B(n816), .C(n815), .Z(n824) );
  IVSVTX4 U1588 ( .A(n1303), .Z(n937) );
  IVSVTX2 U1589 ( .A(n1228), .Z(n1133) );
  ND2SVTX2 U1590 ( .A(n1464), .B(n783), .Z(n750) );
  IVSVTX2 U1591 ( .A(n1005), .Z(n1006) );
  AO17SVTX8 U1592 ( .A(n1706), .B(n1704), .C(n1705), .D(n1773), .Z(n1219) );
  NR3SVTX4 U1593 ( .A(n1134), .B(n1170), .C(n1256), .Z(n744) );
  BFSVTX1 U1594 ( .A(n1560), .Z(n1515) );
  ND2SVTX4 U1595 ( .A(n1486), .B(n1119), .Z(n796) );
  NR2SVTX4 U1596 ( .A(n845), .B(n869), .Z(n726) );
  ND2SVTX4 U1597 ( .A(n1543), .B(n1542), .Z(n1553) );
  ND2SVTX2 U1598 ( .A(n1720), .B(n1119), .Z(n1559) );
  OR2BSVTX4 U1599 ( .A(n1133), .B(n1119), .Z(n1231) );
  CTIVSVTX2 U1600 ( .A(n1140), .Z(n1069) );
  F_AN2SVTX2 U1601 ( .A(n1119), .B(n1493), .Z(n781) );
  IVSVTX2 U1602 ( .A(n1121), .Z(n728) );
  IVSVTX2 U1603 ( .A(n728), .Z(n729) );
  IVSVTX8 U1604 ( .A(n736), .Z(n1321) );
  AO7SVTX4 U1605 ( .A(O[27]), .B(n1588), .C(n1160), .Z(n1161) );
  AO6SVTX8 U1606 ( .A(n756), .B(n1765), .C(n1265), .Z(n1442) );
  F_ND2SVTX0H U1607 ( .A(N[1]), .B(n868), .Z(n980) );
  ND2SVTX4 U1608 ( .A(n1360), .B(n1366), .Z(n1289) );
  IVSVTX6 U1609 ( .A(n1732), .Z(n1733) );
  ND2SVTX2 U1610 ( .A(n1352), .B(n1366), .Z(n1355) );
  AO7SVTX4 U1611 ( .A(n619), .B(n437), .C(n1677), .Z(n1549) );
  CTMUX21NSVTX4 U1612 ( .A(n1108), .B(n1107), .S(n1106), .Z(n1230) );
  ND2SVTX2 U1613 ( .A(n1177), .B(n1313), .Z(n1178) );
  IVSVTX4 U1614 ( .A(n946), .Z(n947) );
  ND3SVTX8 U1615 ( .A(n1345), .B(n1346), .C(n1344), .Z(n1347) );
  ND2SVTX4 U1616 ( .A(n1521), .B(n576), .Z(n1368) );
  AO6ABSVTX8 U1617 ( .A(n1055), .B(n1054), .C(n1053), .Z(n1319) );
  ND2SVTX4 U1618 ( .A(N[8]), .B(n777), .Z(n961) );
  ND2SVTX4 U1619 ( .A(n1648), .B(n1716), .Z(n1649) );
  ND2SVTX4 U1620 ( .A(n1619), .B(n1622), .Z(n735) );
  AO17SVTX6 U1621 ( .A(n782), .B(n1731), .C(n1730), .D(n1729), .Z(n1812) );
  IVSVTX2 U1622 ( .A(n1422), .Z(n757) );
  ND2SVTX2 U1623 ( .A(n1133), .B(n1320), .Z(n1134) );
  CTIVSVTX6 U1624 ( .A(n355), .Z(n950) );
  NR2SVTX2 U1625 ( .A(n1162), .B(n955), .Z(n1163) );
  ND3SVTX8 U1626 ( .A(n725), .B(n911), .C(n946), .Z(n737) );
  IVSVTX4 U1627 ( .A(n1216), .Z(n1162) );
  ND2SVTX4 U1628 ( .A(n1165), .B(n1387), .Z(n1001) );
  AO6SVTX8 U1629 ( .A(n1444), .B(n1693), .C(n1692), .Z(n1503) );
  IVSVTX8 U1630 ( .A(n1428), .Z(n1513) );
  CTBUFSVTX8 U1631 ( .A(n1339), .Z(n974) );
  NR2SVTX2 U1632 ( .A(n1515), .B(n1432), .Z(n1517) );
  ND2SVTX4 U1633 ( .A(n327), .B(n999), .Z(n1165) );
  AO6SVTX2 U1634 ( .A(n1064), .B(n1063), .C(n722), .Z(n1065) );
  ND2SVTX4 U1635 ( .A(n1102), .B(n1101), .Z(n1235) );
  ND3SVTX4 U1636 ( .A(n1233), .B(n1232), .C(n1231), .Z(n1234) );
  IVSVTX2 U1637 ( .A(n1520), .Z(n1316) );
  IVSVTX8 U1638 ( .A(n1323), .Z(n1419) );
  AO7SVTX4 U1639 ( .A(n1525), .B(n1158), .C(n1157), .Z(n1216) );
  IVSVTX2 U1640 ( .A(n1131), .Z(n1132) );
  OR2SVTX2 U1641 ( .A(n1155), .B(n1707), .Z(n1787) );
  IVSVTX0H U1642 ( .A(n1295), .Z(n915) );
  IVSVTX2 U1643 ( .A(n1532), .Z(n1536) );
  IVSVTX4 U1644 ( .A(n1352), .Z(n1334) );
  F_AN2SVTX2 U1645 ( .A(n923), .B(n1294), .Z(n798) );
  NR2SVTX2 U1646 ( .A(n876), .B(n875), .Z(n877) );
  NR2ASVTX2 U1647 ( .A(n1038), .B(n1285), .Z(n886) );
  ND2SVTX2 U1648 ( .A(n1520), .B(n576), .Z(n1353) );
  IVSVTX2 U1649 ( .A(n1391), .Z(n1393) );
  IVSVTX2 U1650 ( .A(n1135), .Z(n740) );
  B_ND2SVTX1 U1651 ( .A(n530), .B(n1613), .Z(n1595) );
  AO6SVTX4 U1652 ( .A(n1727), .B(n1728), .C(n1726), .Z(n1729) );
  F_ND2SVTX1 U1653 ( .A(n1801), .B(n290), .Z(n1807) );
  F_ND2SVTX1 U1654 ( .A(n1797), .B(n1796), .Z(n1799) );
  F_ND2SVTX1 U1655 ( .A(n1698), .B(n1697), .Z(n1700) );
  IVSVTX2 U1656 ( .A(n1742), .Z(n1743) );
  ND3SVTX2 U1657 ( .A(n1540), .B(n1555), .C(n1558), .Z(n1541) );
  NR3ABSVTX8 U1658 ( .A(n1348), .B(n1349), .C(n1347), .Z(n739) );
  NR2SVTX4 U1659 ( .A(n930), .B(n797), .Z(n1305) );
  IVSVTX2 U1660 ( .A(n1036), .Z(n1042) );
  MUX21SVTX4 U1661 ( .A(n1135), .B(n740), .S(n744), .Z(n1136) );
  ND2SVTX4 U1662 ( .A(n282), .B(n272), .Z(n1172) );
  ND2SVTX4 U1663 ( .A(n1413), .B(n1396), .Z(n1377) );
  AN3SVTX4 U1664 ( .A(n1457), .B(n1456), .C(n562), .Z(n783) );
  IVSVTX4 U1665 ( .A(n1495), .Z(n1754) );
  NR2SVTX2 U1666 ( .A(n1454), .B(n1453), .Z(n1457) );
  ND2ASVTX8 U1667 ( .A(n1258), .B(n1098), .Z(n742) );
  ND2ASVTX8 U1668 ( .A(n964), .B(n1294), .Z(n1059) );
  ND2SVTX4 U1669 ( .A(n1294), .B(n1284), .Z(n1333) );
  F_ENSVTX2 U1670 ( .A(n1619), .B(n1627), .Z(n1628) );
  IVSVTX4 U1671 ( .A(n1781), .Z(n1229) );
  AO6SVTX1 U1672 ( .A(N[0]), .B(n943), .C(n1326), .Z(n917) );
  IVSVTX2 U1673 ( .A(n464), .Z(n1514) );
  AO7SVTX4 U1674 ( .A(n1547), .B(n1555), .C(n282), .Z(n1385) );
  ND2SVTX4 U1675 ( .A(n282), .B(n1120), .Z(n1232) );
  ND4ASVTX8 U1676 ( .A(n302), .B(n1232), .C(n1233), .D(n1231), .Z(n1790) );
  ND2SVTX4 U1677 ( .A(n1026), .B(n1027), .Z(n1045) );
  AO7SVTX8 U1678 ( .A(n1562), .B(n1563), .C(n1561), .Z(n1564) );
  NR2SVTX2 U1679 ( .A(n1155), .B(n1707), .Z(n1174) );
  AO7ABSVTX2 U1680 ( .A(n1304), .B(n937), .C(O[28]), .Z(n1308) );
  AO20SVTX4 U1681 ( .A(n1553), .B(n717), .C(n1720), .D(n712), .Z(n1545) );
  AO7SVTX2 U1682 ( .A(n1553), .B(n717), .C(n277), .Z(n1557) );
  AO2ASVTX4 U1683 ( .C(n1366), .D(n962), .A(n1356), .B(n1367), .Z(n1358) );
  ND2SVTX4 U1684 ( .A(n991), .B(n992), .Z(n993) );
  AO4SVTX2 U1685 ( .A(n854), .B(n814), .C(n940), .D(n843), .Z(n815) );
  ND3SVTX4 U1686 ( .A(n922), .B(n924), .C(n832), .Z(n834) );
  AO7NSVTX4 U1687 ( .A(n932), .B(n843), .C(n924), .Z(n925) );
  ND3SVTX8 U1688 ( .A(n807), .B(n806), .C(n805), .Z(n752) );
  AO3NSVTX2 U1689 ( .A(n1329), .B(n1296), .C(n1328), .D(n1327), .Z(n779) );
  IVSVTX4 U1690 ( .A(n1325), .Z(n1329) );
  NR2SVTX2 U1691 ( .A(n1080), .B(n898), .Z(n899) );
  MUX21NSVTX6 U1692 ( .A(n1066), .B(n1065), .S(n1082), .Z(n1250) );
  IVSVTX12 U1693 ( .A(n1073), .Z(n1366) );
  NR2SVTX2 U1694 ( .A(n307), .B(n1070), .Z(n1138) );
  ND2SVTX4 U1695 ( .A(n1145), .B(n541), .Z(n1221) );
  AO7SVTX2 U1696 ( .A(n1012), .B(O[31]), .C(n931), .Z(n934) );
  IVSVTX2 U1697 ( .A(n1320), .Z(n1115) );
  ND2ASVTX8 U1698 ( .A(n1264), .B(n1261), .Z(n756) );
  AO17SVTX8 U1699 ( .A(n1207), .B(n1206), .C(n1205), .D(n1204), .Z(n1704) );
  ND2SVTX2 U1700 ( .A(n1278), .B(n777), .Z(n1282) );
  ND2SVTX2 U1701 ( .A(n1284), .B(n777), .Z(n1288) );
  CTOR3SVTX4 U1702 ( .A(N[5]), .B(N[4]), .C(n1031), .Z(n778) );
  ND2SVTX4 U1703 ( .A(n1034), .B(n1000), .Z(n1121) );
  F_ND2SVTX1 U1704 ( .A(n1780), .B(n1781), .Z(n1786) );
  ND3SVTX4 U1705 ( .A(n1718), .B(n753), .C(n764), .Z(n1605) );
  ND2ASVTX8 U1706 ( .A(n758), .B(n1240), .Z(n1444) );
  IVSVTX4 U1707 ( .A(n863), .Z(n759) );
  BFSVTX1 U1708 ( .A(n1625), .Z(n1593) );
  AO6SVTX2 U1709 ( .A(n1593), .B(n1592), .C(n711), .Z(n1594) );
  AO6SVTX2 U1710 ( .A(n1615), .B(n1625), .C(n1614), .Z(n1616) );
  OR3SVTX4 U1711 ( .A(n1274), .B(n1072), .C(n934), .Z(n762) );
  NR2SVTX2 U1712 ( .A(n998), .B(n754), .Z(n999) );
  NR2SVTX4 U1713 ( .A(n909), .B(n983), .Z(n946) );
  NR2ASVTX6 U1714 ( .A(n1367), .B(n1299), .Z(n1392) );
  IVSVTX4 U1715 ( .A(n1161), .Z(n1540) );
  IVSVTX6 U1716 ( .A(n1540), .Z(n1617) );
  AO6NSVTX1 U1717 ( .A(n1706), .B(n1802), .C(n1705), .Z(n1788) );
  AO6SVTX1 U1718 ( .A(n1788), .B(n1775), .C(n1774), .Z(n1776) );
  ND2SVTX2 U1719 ( .A(n1026), .B(n1027), .Z(n1028) );
  AO7SVTX1 U1720 ( .A(n1805), .B(n1804), .C(n1803), .Z(n1806) );
  NR2SVTX2 U1721 ( .A(n970), .B(n586), .Z(n930) );
  ND2SVTX2 U1722 ( .A(n981), .B(n587), .Z(n874) );
  NR2SVTX2 U1723 ( .A(n1808), .B(n1459), .Z(n1462) );
  ND3ABSVTX4 U1724 ( .A(n895), .B(n893), .C(n307), .Z(n897) );
  F_ND2SVTX1 U1725 ( .A(n1769), .B(n1768), .Z(n1771) );
  ND2SVTX2 U1726 ( .A(n1567), .B(n1622), .Z(n1568) );
  FAS1SVTX4 U1727 ( .A(n1677), .B(n755), .CI(n1675), .CO(n1719), .Z(n1674) );
  ND2SVTX2 U1728 ( .A(n1428), .B(n1119), .Z(n1423) );
  NR2SVTX2 U1729 ( .A(n942), .B(n903), .Z(n905) );
  ND2SVTX4 U1730 ( .A(n1285), .B(n763), .Z(n903) );
  AO7SVTX8 U1731 ( .A(n1443), .B(n1442), .C(n1441), .Z(n1692) );
  F_ND2SVTX1 U1732 ( .A(n1691), .B(n1690), .Z(n1696) );
  NR2SVTX2 U1733 ( .A(n307), .B(n1446), .Z(n1125) );
  IVSVTX4 U1734 ( .A(n1033), .Z(n1446) );
  ND2SVTX4 U1735 ( .A(n1111), .B(n1052), .Z(n1228) );
  EOSVTX8 U1736 ( .A(n1814), .B(n1813), .Z(O[26]) );
  ND3ABSVTX4 U1737 ( .A(n327), .B(n1071), .C(n896), .Z(n1150) );
  NR3SVTX2 U1738 ( .A(n1314), .B(O[29]), .C(n1315), .Z(n1309) );
  ND2SVTX4 U1739 ( .A(n1499), .B(n1498), .Z(n1750) );
  IVSVTX2 U1740 ( .A(n892), .Z(n893) );
  IVSVTX2 U1741 ( .A(n1618), .Z(n1639) );
  ND2SVTX2 U1742 ( .A(n1747), .B(n1746), .Z(n1748) );
  ND2SVTX2 U1743 ( .A(n1119), .B(n1609), .Z(n1422) );
  ND2SVTX2 U1744 ( .A(n1603), .B(n1119), .Z(n1383) );
  ND2SVTX2 U1745 ( .A(n1150), .B(n1140), .Z(n1151) );
  BFSVTX2 U1746 ( .A(N[18]), .Z(n963) );
  AN2SVTX0H U1747 ( .A(n1606), .B(n1724), .Z(n780) );
  AN2SVTX4 U1748 ( .A(n1220), .B(n1119), .Z(n792) );
  OR2SVTX1 U1749 ( .A(n312), .B(n964), .Z(n793) );
  AO7SVTX2 U1750 ( .A(n929), .B(O[31]), .C(n928), .Z(n797) );
  IVSVTX2 U1751 ( .A(n1361), .Z(n969) );
  F_AN2SVTX2 U1752 ( .A(n1020), .B(n1285), .Z(n802) );
  NR2SVTX6 U1753 ( .A(n675), .B(n870), .Z(n806) );
  ND2ASVTX8 U1754 ( .A(N[25]), .B(n804), .Z(n869) );
  IVSVTX6 U1755 ( .A(N[10]), .Z(n964) );
  NR2SVTX8 U1756 ( .A(N[9]), .B(N[11]), .Z(n810) );
  NR2SVTX4 U1757 ( .A(N[7]), .B(N[6]), .Z(n827) );
  NR2SVTX4 U1758 ( .A(N[5]), .B(N[4]), .Z(n828) );
  NR2SVTX4 U1759 ( .A(N[15]), .B(N[14]), .Z(n813) );
  ND2SVTX4 U1760 ( .A(n813), .B(n881), .Z(n854) );
  BFSVTX6 U1761 ( .A(N[9]), .Z(n972) );
  ND2SVTX4 U1762 ( .A(n312), .B(n819), .Z(n991) );
  AO6CSVTX8 U1763 ( .A(n312), .B(n821), .C(n820), .Z(n992) );
  BFSVTX2 U1764 ( .A(N[17]), .Z(n927) );
  ND2SVTX2 U1765 ( .A(n927), .B(n861), .Z(n823) );
  IVSVTX4 U1766 ( .A(n1277), .Z(n825) );
  AN2SVTX8 U1767 ( .A(n828), .B(n827), .Z(n857) );
  NR2SVTX4 U1768 ( .A(n834), .B(n833), .Z(n835) );
  IVSVTX4 U1769 ( .A(N[23]), .Z(n931) );
  IVSVTX4 U1770 ( .A(n931), .Z(n1314) );
  ND2SVTX4 U1771 ( .A(n840), .B(n839), .Z(n841) );
  IVSVTX4 U1772 ( .A(N[13]), .Z(n843) );
  ND3SVTX6 U1773 ( .A(N[11]), .B(n843), .C(n808), .Z(n844) );
  AO7SVTX6 U1774 ( .A(n856), .B(n857), .C(n855), .Z(n858) );
  BFSVTX2 U1775 ( .A(N[10]), .Z(n882) );
  IVSVTX2 U1776 ( .A(n1059), .Z(n876) );
  ND2SVTX2 U1777 ( .A(n940), .B(n1294), .Z(n1063) );
  AN2SVTX4 U1778 ( .A(n1064), .B(n1063), .Z(n1361) );
  AO6SVTX2 U1779 ( .A(n882), .B(n881), .C(n940), .Z(n883) );
  NR2SVTX8 U1780 ( .A(n754), .B(n945), .Z(n949) );
  BFSVTX6 U1781 ( .A(N[11]), .Z(n1278) );
  IVSVTX4 U1782 ( .A(n1047), .Z(n889) );
  ND3SVTX6 U1783 ( .A(n307), .B(n1139), .C(n1124), .Z(n890) );
  ND2SVTX4 U1784 ( .A(n1014), .B(n1015), .Z(n1034) );
  ND2SVTX4 U1785 ( .A(n899), .B(n900), .Z(n1258) );
  AO7SVTX2 U1786 ( .A(n941), .B(n1325), .C(n705), .Z(n906) );
  NR2ASVTX4 U1787 ( .A(n720), .B(n1291), .Z(n904) );
  BFSVTX1 U1788 ( .A(N[20]), .Z(n1295) );
  IVSVTX4 U1789 ( .A(n952), .Z(n926) );
  IVSVTX4 U1790 ( .A(n803), .Z(n936) );
  ND2SVTX4 U1791 ( .A(n1304), .B(n937), .Z(n938) );
  ND2ASVTX8 U1792 ( .A(n722), .B(n948), .Z(n1356) );
  NR2SVTX8 U1793 ( .A(n1590), .B(n951), .Z(n1097) );
  ND2SVTX2 U1794 ( .A(n963), .B(n1294), .Z(n967) );
  ND2SVTX4 U1795 ( .A(n1370), .B(n1522), .Z(n976) );
  IVSVTX4 U1796 ( .A(n992), .Z(n984) );
  NR2ASVTX1 U1797 ( .A(N[4]), .B(n312), .Z(n989) );
  ND2SVTX2 U1798 ( .A(N[3]), .B(n1294), .Z(n998) );
  IVSVTX4 U1799 ( .A(n1009), .Z(n1276) );
  ND2SVTX8 U1800 ( .A(n1008), .B(n1007), .Z(n1181) );
  NR2SVTX8 U1801 ( .A(n1181), .B(n1011), .Z(n1091) );
  MUX21NSVTX6 U1802 ( .A(n1023), .B(n1013), .S(n1043), .Z(n1156) );
  AO7ABSVTX2 U1803 ( .A(n484), .B(n1326), .C(n1017), .Z(n1026) );
  ND2SVTX6 U1804 ( .A(n1025), .B(n1024), .Z(n1044) );
  IVSVTX2 U1805 ( .A(n1046), .Z(n1041) );
  ND3ABSVTX8 U1806 ( .A(n1057), .B(n1056), .C(n1319), .Z(n1255) );
  IVSVTX2 U1807 ( .A(n1076), .Z(n1060) );
  NR3SVTX8 U1808 ( .A(n1080), .B(n1078), .C(n1079), .Z(n1087) );
  EOSVTX8 U1809 ( .A(n1493), .B(n1090), .Z(n1473) );
  ND2ASVTX8 U1810 ( .A(n1468), .B(n1092), .Z(n1476) );
  ND2SVTX6 U1811 ( .A(n1104), .B(n1103), .Z(n1113) );
  ND2SVTX4 U1812 ( .A(n1483), .B(n1136), .Z(n1233) );
  ND4ABSVTX8 U1813 ( .A(n1225), .B(n1228), .C(n1224), .D(n1226), .Z(n1781) );
  NR2SVTX4 U1814 ( .A(n1800), .B(n1805), .Z(n1706) );
  ND3ABSVTX4 U1815 ( .A(n955), .B(n1161), .C(n1201), .Z(n1195) );
  IVSVTX4 U1816 ( .A(n1772), .Z(n1217) );
  ND2SVTX4 U1817 ( .A(n1236), .B(n1790), .Z(n1237) );
  NR2SVTX2 U1818 ( .A(n1248), .B(n1247), .Z(n1253) );
  ENSVTX8 U1819 ( .A(n1486), .B(n1257), .Z(n1269) );
  ND2SVTX6 U1820 ( .A(n1769), .B(n756), .Z(n1434) );
  ND2ASVTX8 U1821 ( .A(n1135), .B(n1263), .Z(n1768) );
  IVSVTX8 U1822 ( .A(n1764), .Z(n1265) );
  ND2SVTX4 U1823 ( .A(n674), .B(n802), .Z(n1286) );
  ND2SVTX2 U1824 ( .A(n1295), .B(n1294), .Z(n1327) );
  ND2ASVTX8 U1825 ( .A(n1297), .B(n791), .Z(n1364) );
  AO2SVTX2 U1826 ( .A(n748), .B(n1364), .C(n1520), .D(n1371), .Z(n1530) );
  AO2SVTX2 U1827 ( .A(n1522), .B(n1300), .C(n1366), .D(n1521), .Z(n1302) );
  B_ND2SVTX2 U1828 ( .A(n1523), .B(n471), .Z(n1301) );
  IVSVTX4 U1829 ( .A(n1364), .Z(n1357) );
  ND2ASVTX8 U1830 ( .A(n1533), .B(n1318), .Z(n1603) );
  ND2SVTX4 U1831 ( .A(n1320), .B(n1319), .Z(n1400) );
  ND2SVTX4 U1832 ( .A(n1360), .B(n576), .Z(n1406) );
  NR2SVTX4 U1833 ( .A(n212), .B(n1405), .Z(n1338) );
  ND2ASVTX8 U1834 ( .A(n1336), .B(n624), .Z(n1408) );
  ND4ABSVTX8 U1835 ( .A(n1400), .B(n1466), .C(n1419), .D(n1417), .Z(n1350) );
  ND2SVTX4 U1836 ( .A(n1360), .B(n1522), .Z(n1354) );
  ND2SVTX4 U1837 ( .A(n1360), .B(n1371), .Z(n1391) );
  ND2SVTX4 U1838 ( .A(n1391), .B(n1390), .Z(n1375) );
  ND2SVTX4 U1839 ( .A(n1371), .B(n1370), .Z(n1362) );
  ND2SVTX4 U1840 ( .A(n962), .B(n1371), .Z(n1372) );
  NR2SVTX4 U1841 ( .A(n1411), .B(n1394), .Z(n1373) );
  ND3ABSVTX8 U1842 ( .A(n1379), .B(n1380), .C(n785), .Z(n1381) );
  NR2SVTX6 U1843 ( .A(n1400), .B(n1466), .Z(n1418) );
  ND2SVTX4 U1844 ( .A(n1555), .B(n1542), .Z(n1401) );
  NR2SVTX4 U1845 ( .A(n1449), .B(n1413), .Z(n1409) );
  ND2ASVTX8 U1846 ( .A(n1411), .B(n1410), .Z(n1609) );
  IVSVTX4 U1847 ( .A(n1609), .Z(n1451) );
  ND2SVTX4 U1848 ( .A(n1431), .B(n1430), .Z(n1509) );
  ND2SVTX4 U1849 ( .A(n742), .B(n1437), .Z(n1433) );
  NR2SVTX8 U1850 ( .A(n1434), .B(n1433), .Z(n1693) );
  AO6SVTX8 U1851 ( .A(n702), .B(n1440), .C(n1439), .Z(n1441) );
  NR2SVTX4 U1852 ( .A(n1445), .B(n1447), .Z(n1454) );
  ND2ASVTX8 U1853 ( .A(n1496), .B(n1754), .Z(n1463) );
  ENSVTX8 U1854 ( .A(n1472), .B(n1471), .Z(n1477) );
  ND2ASVTX8 U1855 ( .A(n278), .B(n1477), .Z(n1489) );
  IVSVTX2 U1856 ( .A(n1492), .Z(n1691) );
  ND2SVTX4 U1857 ( .A(n1698), .B(n1691), .Z(n1751) );
  IVSVTX4 U1858 ( .A(n1751), .Z(n1485) );
  ND2SVTX6 U1859 ( .A(n273), .B(n1485), .Z(n1502) );
  ND2SVTX4 U1860 ( .A(n1609), .B(n1608), .Z(n1510) );
  ND3SVTX2 U1861 ( .A(n1529), .B(n1530), .C(n1531), .Z(n1538) );
  NR2SVTX4 U1862 ( .A(n1534), .B(n1533), .Z(n1535) );
  ND2SVTX4 U1863 ( .A(n1543), .B(n279), .Z(n1539) );
  IVSVTX4 U1864 ( .A(n1539), .Z(n1558) );
  NR2SVTX4 U1865 ( .A(n437), .B(n1541), .Z(n1676) );
  NR2SVTX4 U1866 ( .A(n279), .B(n1575), .Z(n1567) );
  IVSVTX4 U1867 ( .A(n1553), .Z(n1554) );
  AO6SVTX8 U1868 ( .A(n1565), .B(n1570), .C(n1564), .Z(n1623) );
  ND2ASVTX8 U1869 ( .A(n1575), .B(n1620), .Z(n1576) );
  IVSVTX2 U1870 ( .A(n1575), .Z(n1619) );
  ENSVTX8 U1871 ( .A(n277), .B(n1578), .Z(n1646) );
  IVSVTX2 U1872 ( .A(n1645), .Z(n1597) );
  ND2SVTX2 U1873 ( .A(n1597), .B(n1643), .Z(n1598) );
  ENSVTX4 U1874 ( .A(n403), .B(n1598), .Z(O[18]) );
  NR2ASVTX8 U1875 ( .A(n1667), .B(n1666), .Z(n1669) );
  AO6CSVTX4 U1876 ( .A(n1741), .B(n320), .C(n708), .Z(n1671) );
  EOSVTX8 U1877 ( .A(n1672), .B(n1671), .Z(O[22]) );
  AO6SVTX4 U1878 ( .A(n1741), .B(n1686), .C(n1685), .Z(n1687) );
  EOSVTX8 U1879 ( .A(n1688), .B(n1687), .Z(O[24]) );
  AO6SVTX1 U1880 ( .A(n1770), .B(n1693), .C(n1692), .Z(n1699) );
  NR2SVTX6 U1881 ( .A(n1725), .B(n1722), .Z(n1728) );
  AO7SVTX4 U1882 ( .A(n1725), .B(n1724), .C(n1723), .Z(n1726) );
  ENSVTX4 U1883 ( .A(n794), .B(n1812), .Z(O[25]) );
  IVSVTX2 U1884 ( .A(n1734), .Z(n1744) );
  AO7SVTX2 U1885 ( .A(n1744), .B(n732), .C(n1736), .Z(n1737) );
  ENSVTX4 U1886 ( .A(n1738), .B(n1737), .Z(O[20]) );
  ND2SVTX2 U1887 ( .A(n708), .B(n320), .Z(n1740) );
  ENSVTX4 U1888 ( .A(n1741), .B(n1740), .Z(O[21]) );
  EOSVTX4 U1889 ( .A(n1744), .B(n1743), .Z(O[19]) );
  F_ND2SVTX1 U1890 ( .A(n1749), .B(n1750), .Z(n1758) );
  F_ND2SVTX1 U1891 ( .A(n238), .B(n1764), .Z(n1767) );
endmodule

