
module remap_top ( num_i, rslt_o );
  input [31:0] num_i;
  output [31:0] rslt_o;
  wire   n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n428, n429, n430,
         n431, n432, n433, n434, n438, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n450, n451, n452, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n749, n750, n751, n752, n753, n754, n755, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n814, n815, n816, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n856, n857, n859, n860, n861, n862, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n894, n895, n896, n898, n899, n900, n902,
         n903, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n930, n931, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1092, n1093, n1094, n1095, n1096,
         n1097, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1453, n1454, n1455, n1456, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1918, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1953, n1954, n1955, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307;

  BFSVTX0H U417 ( .A(n2636), .Z(rslt_o[29]) );
  AO7SVTX4 U418 ( .A(n4188), .B(n4187), .C(n4186), .Z(rslt_o[26]) );
  B_ND2SVTX2 U419 ( .A(n4201), .B(n4200), .Z(n4202) );
  IVSVTX1 U420 ( .A(n4203), .Z(n4212) );
  B_ND2SVTX2 U421 ( .A(n450), .B(n4266), .Z(n4267) );
  IVSVTX0H U422 ( .A(n4262), .Z(n4263) );
  IVSVTX2 U423 ( .A(n1873), .Z(n2432) );
  IVSVTX2 U424 ( .A(n339), .Z(n4304) );
  IVSVTX2 U425 ( .A(n2376), .Z(n4201) );
  IVSVTX0H U426 ( .A(n4305), .Z(n4285) );
  F_ND2ASVTX2 U427 ( .A(n1350), .B(n1351), .Z(n4200) );
  IVSVTX0H U428 ( .A(n4254), .Z(n4251) );
  IVSVTX0H U429 ( .A(n4297), .Z(n4298) );
  IVSVTX0H U430 ( .A(n4288), .Z(n1250) );
  NR2ASVTX2 U431 ( .A(n1350), .B(n1351), .Z(n2376) );
  ND2SVTX4 U432 ( .A(n1456), .B(n1451), .Z(n3109) );
  ND2SVTX2 U433 ( .A(n4067), .B(n392), .Z(n4189) );
  BFSVTX2 U434 ( .A(n1716), .Z(n413) );
  ND2ASVTX4 U435 ( .A(n763), .B(n953), .Z(n4283) );
  NR2ASVTX1 U436 ( .A(n514), .B(n3260), .Z(n4168) );
  AN3SVTX2 U437 ( .A(n1715), .B(n4096), .C(n4167), .Z(n490) );
  NR2ASVTX1 U438 ( .A(n506), .B(n3147), .Z(n4146) );
  NR2ASVTX4 U439 ( .A(n4051), .B(n1582), .Z(n1464) );
  NR2ASVTX4 U440 ( .A(n763), .B(n953), .Z(n4281) );
  B_ND2SVTX2 U441 ( .A(n2212), .B(n2213), .Z(n368) );
  IVSVTX0H U442 ( .A(n4180), .Z(n2303) );
  F_AN2SVTX2 U443 ( .A(n4098), .B(n4097), .Z(n1746) );
  ND3SVTX4 U444 ( .A(n1445), .B(n2005), .C(n2002), .Z(n1444) );
  AN2SVTX2 U445 ( .A(n506), .B(n4128), .Z(n498) );
  ND2SVTX1 U446 ( .A(n4066), .B(n4065), .Z(n1704) );
  AO6SVTX6 U447 ( .A(n1668), .B(n4294), .C(n1891), .Z(n2434) );
  ND2ASVTX4 U448 ( .A(n2195), .B(n2194), .Z(n3200) );
  NR2ASVTX1 U449 ( .A(n1422), .B(n4160), .Z(n4156) );
  IVSVTX2 U450 ( .A(n1304), .Z(n2194) );
  IVSVTX2 U451 ( .A(n4078), .Z(n4081) );
  NR2ASVTX1 U452 ( .A(n4174), .B(n4093), .Z(n4094) );
  AO7CNSVTX4 U453 ( .A(n622), .B(n3145), .C(n1660), .Z(n2213) );
  ND3SVTX1 U454 ( .A(n4174), .B(n2349), .C(n1715), .Z(n4097) );
  IVSVTX0H U455 ( .A(n4172), .Z(n4098) );
  B_ND2SVTX2 U456 ( .A(n4142), .B(n4144), .Z(n1445) );
  ND2SVTX2 U457 ( .A(n642), .B(n3298), .Z(n1628) );
  IVSVTX0H U458 ( .A(n4135), .Z(n2159) );
  ND3SVTX6 U459 ( .A(n4230), .B(n4235), .C(n2102), .Z(n3717) );
  NR2ASVTX2 U460 ( .A(n4176), .B(n4115), .Z(n4180) );
  NR2ASVTX1 U461 ( .A(n2248), .B(n3528), .Z(n764) );
  NR2ASVTX2 U462 ( .A(n4174), .B(n3260), .Z(n4096) );
  AO6CSVTX6 U463 ( .A(n1408), .B(n1404), .C(n529), .Z(n1407) );
  NR2SVTX2 U464 ( .A(n1660), .B(n4130), .Z(n1783) );
  CTBUFSVTX2 U465 ( .A(n1596), .Z(n367) );
  AO7SVTX4 U466 ( .A(n3262), .B(n3263), .C(n2214), .Z(n937) );
  AO7SVTX2 U467 ( .A(n4059), .B(n1641), .C(n1899), .Z(n2219) );
  ND3SVTX1 U468 ( .A(n4163), .B(n4160), .C(n3132), .Z(n1911) );
  AO7SVTX2 U469 ( .A(n3108), .B(n525), .C(n3106), .Z(n1454) );
  AO7SVTX4 U470 ( .A(n1929), .B(n1927), .C(n392), .Z(n1926) );
  IVSVTX2 U471 ( .A(n2103), .Z(n1350) );
  NR2SVTX2 U472 ( .A(n3260), .B(n3297), .Z(n3298) );
  AO7SVTX2 U473 ( .A(n4154), .B(n4153), .C(n4152), .Z(n4162) );
  ND2ASVTX4 U474 ( .A(n523), .B(n3164), .Z(n4078) );
  ND2SVTX2 U475 ( .A(n4167), .B(n454), .Z(n784) );
  F_IVSVTX1 U476 ( .A(n1705), .Z(n4093) );
  IVSVTX0H U477 ( .A(n3351), .Z(n3213) );
  IVSVTX2 U478 ( .A(n3108), .Z(n1646) );
  CTIVSVTX2 U479 ( .A(n3163), .Z(n1460) );
  CTIVSVTX2 U480 ( .A(n1637), .Z(n1927) );
  IVSVTX0H U481 ( .A(n1494), .Z(n571) );
  ND2SVTX2 U482 ( .A(n3293), .B(n2453), .Z(n3295) );
  ND2SVTX2 U483 ( .A(n3057), .B(n3179), .Z(n889) );
  NR3ABSVTX6 U484 ( .A(n3113), .B(n2053), .C(n1462), .Z(n2210) );
  ND3SVTX2 U485 ( .A(n1590), .B(n558), .C(n1589), .Z(n2182) );
  AO7SVTX4 U486 ( .A(n2349), .B(n4069), .C(n497), .Z(n1408) );
  NR2SVTX2 U487 ( .A(n615), .B(n4125), .Z(n4130) );
  AN3SVTX1 U488 ( .A(n530), .B(n3278), .C(n3277), .Z(n3296) );
  NR3ABSVTX4 U489 ( .A(n1013), .B(n2445), .C(n1011), .Z(n1009) );
  NR4ABSVTX4 U490 ( .A(n4171), .B(n3410), .C(n4167), .D(n1843), .Z(n375) );
  ND2ASVTX4 U491 ( .A(n3260), .B(n3164), .Z(n4077) );
  AN2SVTX2 U492 ( .A(n3305), .B(n3367), .Z(n3309) );
  BFSVTX2 U493 ( .A(n2362), .Z(n401) );
  NR2SVTX2 U494 ( .A(n4108), .B(n4153), .Z(n1574) );
  AO3SVTX2 U495 ( .A(n4104), .B(n1270), .C(n4103), .D(n4102), .Z(n1929) );
  NR3ABSVTX2 U496 ( .A(n3057), .B(n3106), .C(n560), .Z(n3107) );
  ND2ASVTX6 U497 ( .A(n523), .B(n2400), .Z(n3120) );
  IVSVTX0H U498 ( .A(n4092), .Z(n1589) );
  IVSVTX2 U499 ( .A(n3331), .Z(n789) );
  BFSVTX2 U500 ( .A(n2291), .Z(n1660) );
  IVSVTX2 U501 ( .A(n2055), .Z(n1462) );
  F_ND3SVTX2 U502 ( .A(n1928), .B(n4105), .C(n4058), .Z(n1637) );
  IVSVTX0H U503 ( .A(n4163), .Z(n594) );
  IVSVTX0H U504 ( .A(n4108), .Z(n1931) );
  NR2SVTX4 U505 ( .A(n3163), .B(n2134), .Z(n4085) );
  IVSVTX4 U506 ( .A(n3972), .Z(n566) );
  NR2SVTX2 U507 ( .A(n4140), .B(n4139), .Z(n1175) );
  NR3SVTX6 U508 ( .A(n1846), .B(n1847), .C(n3408), .Z(n1844) );
  ND2SVTX2 U509 ( .A(n977), .B(n489), .Z(n982) );
  ND3SVTX4 U510 ( .A(n2438), .B(n976), .C(n975), .Z(n979) );
  ND3SVTX4 U511 ( .A(n523), .B(n1734), .C(n3299), .Z(n1733) );
  CTIVSVTX2 U512 ( .A(n4079), .Z(n3113) );
  BFSVTX2 U513 ( .A(n2061), .Z(n1172) );
  ND3SVTX6 U514 ( .A(n1899), .B(n1161), .C(n1160), .Z(n1159) );
  NR2SVTX2 U515 ( .A(n1635), .B(n4175), .Z(n4110) );
  IVSVTX4 U516 ( .A(n4257), .Z(n2367) );
  AO7CSVTX4 U517 ( .A(n3342), .B(n741), .C(n3387), .Z(n2453) );
  BFSVTX2 U518 ( .A(n4057), .Z(n1641) );
  ND3SVTX2 U519 ( .A(n3275), .B(n3274), .C(n1932), .Z(n3278) );
  NR2SVTX4 U520 ( .A(n4107), .B(n4159), .Z(n3108) );
  IVSVTX0H U521 ( .A(n4150), .Z(n4154) );
  NR2SVTX2 U522 ( .A(n1588), .B(n573), .Z(n1590) );
  NR2ASVTX2 U523 ( .A(n4116), .B(n4115), .Z(n4126) );
  ND2ASVTX4 U524 ( .A(n2233), .B(n1694), .Z(n3761) );
  ND4ASVTX4 U525 ( .A(n1466), .B(n2084), .C(n1282), .D(n1281), .Z(n1280) );
  ND4ABSVTX6 U526 ( .A(n1833), .B(n3688), .C(n1832), .D(n1831), .Z(n1946) );
  AO6SVTX2 U527 ( .A(n2236), .B(n530), .C(n3389), .Z(n2235) );
  BFSVTX2 U528 ( .A(n2083), .Z(n392) );
  ND2ASVTX1 U529 ( .A(n1932), .B(n2103), .Z(n2433) );
  ND2SVTX4 U530 ( .A(n3528), .B(n1084), .Z(n797) );
  IVSVTX2 U531 ( .A(n4174), .Z(n579) );
  NR2ASVTX1 U532 ( .A(n3342), .B(n1932), .Z(n3276) );
  NR2SVTX2 U533 ( .A(n1531), .B(n3528), .Z(n2386) );
  NR2SVTX2 U534 ( .A(n3377), .B(n509), .Z(n1862) );
  NR2ASVTX1 U535 ( .A(n506), .B(n4120), .Z(n4176) );
  ND2ASVTX6 U536 ( .A(n534), .B(n4151), .Z(n4107) );
  IVSVTX6 U537 ( .A(n1461), .Z(n4091) );
  CTIVSVTX2 U538 ( .A(n1246), .Z(n4063) );
  IVSVTX2 U539 ( .A(n3347), .Z(n529) );
  IVSVTX2 U540 ( .A(n3316), .Z(n883) );
  CTIVSVTX2 U541 ( .A(n3193), .Z(n3194) );
  CTIVSVTX2 U542 ( .A(n3307), .Z(n3305) );
  IVSVTX6 U543 ( .A(n642), .Z(n1896) );
  CTIVSVTX2 U544 ( .A(n3294), .Z(n3259) );
  IVSVTX0H U545 ( .A(n3342), .Z(n3274) );
  IVSVTX0H U546 ( .A(n4057), .Z(n3222) );
  IVSVTX0H U547 ( .A(n4041), .Z(n4038) );
  ND2SVTX2 U548 ( .A(n4055), .B(n4056), .Z(n4059) );
  ND2SVTX2 U549 ( .A(n2248), .B(n3972), .Z(n4048) );
  IVSVTX2 U550 ( .A(n2023), .Z(n870) );
  ND2SVTX2 U551 ( .A(n4135), .B(n4174), .Z(n3019) );
  ND3ABSVTX6 U552 ( .A(n4139), .B(n2932), .C(n1245), .Z(n1160) );
  ND2ASVTX4 U553 ( .A(n1676), .B(n3948), .Z(n1158) );
  ND2SVTX4 U554 ( .A(n3907), .B(n3561), .Z(n4250) );
  IVSVTX0H U555 ( .A(n3341), .Z(n3275) );
  ND3SVTX2 U556 ( .A(n3344), .B(n3343), .C(n3345), .Z(n791) );
  IVSVTX4 U557 ( .A(n1557), .Z(n1554) );
  NR2SVTX6 U558 ( .A(n3528), .B(n1084), .Z(n4262) );
  F_ND2SVTX0H U559 ( .A(n564), .B(n1264), .Z(n3236) );
  IVSVTX4 U560 ( .A(n3143), .Z(n4115) );
  ND2SVTX2 U561 ( .A(n3141), .B(n1255), .Z(n2084) );
  ND2ASVTX4 U562 ( .A(n509), .B(n3013), .Z(n4109) );
  ND2SVTX2 U563 ( .A(n3330), .B(n3328), .Z(n3329) );
  ND4SVTX4 U564 ( .A(n3777), .B(n3778), .C(n3776), .D(n3775), .Z(n3807) );
  AO6SVTX6 U565 ( .A(n2349), .B(n1705), .C(n4069), .Z(n3348) );
  AN3SVTX4 U566 ( .A(n1328), .B(n793), .C(n3117), .Z(n2361) );
  AO6ASVTX6 U567 ( .A(n2363), .B(n3727), .C(n2382), .Z(n3734) );
  AO7ABSVTX2 U568 ( .A(n3311), .B(n2352), .C(n3346), .Z(n792) );
  NR3ABSVTX4 U569 ( .A(n1494), .B(n1705), .C(n2056), .Z(n2400) );
  ND2SVTX2 U570 ( .A(n2276), .B(n565), .Z(n3350) );
  F_AN2SVTX2 U571 ( .A(n3111), .B(n3112), .Z(n4079) );
  ND2SVTX2 U572 ( .A(n3312), .B(n1303), .Z(n3315) );
  NR2SVTX2 U573 ( .A(n3133), .B(n1276), .Z(n1275) );
  ND3SVTX4 U574 ( .A(n2026), .B(n3335), .C(n4159), .Z(n2022) );
  B_ND2SVTX2 U575 ( .A(n350), .B(n3354), .Z(n837) );
  AO6CSVTX4 U576 ( .A(n1603), .B(n3379), .C(n1602), .Z(n2438) );
  ND3ABSVTX4 U577 ( .A(n3254), .B(n3251), .C(n1235), .Z(n3256) );
  ND3ABSVTX4 U578 ( .A(n3381), .B(n524), .C(n3303), .Z(n975) );
  AO6NSVTX4 U579 ( .A(n2054), .B(n2378), .C(n4070), .Z(n466) );
  IVSVTX4 U580 ( .A(n524), .Z(n1899) );
  IVSVTX2 U581 ( .A(n793), .Z(n2113) );
  CTIVSVTX2 U582 ( .A(n2932), .Z(n572) );
  IVSVTX6 U583 ( .A(n1597), .Z(n2346) );
  IVSVTX2 U584 ( .A(n3688), .Z(n522) );
  ND2ASVTX6 U585 ( .A(n1866), .B(n647), .Z(n1874) );
  IVSVTX2 U586 ( .A(n509), .Z(n2167) );
  IVSVTX2 U587 ( .A(n3407), .Z(n3397) );
  CTIVSVTX2 U588 ( .A(n3185), .Z(n3186) );
  IVSVTX2 U589 ( .A(n2101), .Z(n1833) );
  IVSVTX2 U590 ( .A(n2426), .Z(n1603) );
  IVSVTX2 U591 ( .A(n2058), .Z(n3115) );
  IVSVTX0H U592 ( .A(n4055), .Z(n1288) );
  IVSVTX2 U593 ( .A(n1532), .Z(n1531) );
  IVSVTX2 U594 ( .A(n2252), .Z(n717) );
  IVSVTX2 U595 ( .A(n3168), .Z(n4105) );
  NR2ASVTX4 U596 ( .A(n596), .B(n3369), .Z(n3316) );
  NR2SVTX4 U597 ( .A(n3321), .B(n573), .Z(n3347) );
  NR2SVTX2 U598 ( .A(n2027), .B(n3333), .Z(n2026) );
  NR2SVTX2 U599 ( .A(n3223), .B(n580), .Z(n3239) );
  ND3SVTX6 U600 ( .A(n2429), .B(n3921), .C(n3922), .Z(n397) );
  ND2SVTX2 U601 ( .A(n793), .B(n3948), .Z(n2114) );
  AO6SVTX6 U602 ( .A(n3735), .B(n3736), .C(n2382), .Z(n3760) );
  B_ND2SVTX2 U603 ( .A(n464), .B(n3936), .Z(n905) );
  NR2ASVTX4 U604 ( .A(n2932), .B(n4141), .Z(n1162) );
  B_ND2SVTX2 U605 ( .A(n735), .B(n3985), .Z(n3992) );
  ND2SVTX2 U606 ( .A(n712), .B(n711), .Z(n3579) );
  AN2SVTX4 U607 ( .A(n4066), .B(n3990), .Z(n2441) );
  NR2ASVTX6 U608 ( .A(n507), .B(n3112), .Z(n4092) );
  AN3SVTX4 U609 ( .A(n3878), .B(n3879), .C(n1864), .Z(n493) );
  IVSVTX4 U610 ( .A(n1953), .Z(n3528) );
  AN2SVTX4 U611 ( .A(n4022), .B(n3845), .Z(n1461) );
  B_ND2SVTX2 U612 ( .A(n910), .B(n1235), .Z(n3252) );
  AO6SVTX4 U613 ( .A(n3770), .B(n3773), .C(n524), .Z(n3777) );
  CTBUFSVTX2 U614 ( .A(n2936), .Z(n445) );
  NR2SVTX2 U615 ( .A(n1293), .B(n3353), .Z(n350) );
  IVSVTX2 U616 ( .A(n477), .Z(n1289) );
  ND3ABSVTX6 U617 ( .A(n2136), .B(n1910), .C(n3845), .Z(n2135) );
  BFSVTX2 U618 ( .A(n3739), .Z(n865) );
  BFSVTX8 U619 ( .A(n2067), .Z(n733) );
  AO6CSVTX4 U620 ( .A(n1864), .B(n3929), .C(n3793), .Z(n2105) );
  IVSVTX8 U621 ( .A(n2350), .Z(n523) );
  IVSVTX2 U622 ( .A(n3165), .Z(n532) );
  IVSVTX0H U623 ( .A(n622), .Z(n1560) );
  IVSVTX2 U624 ( .A(n2250), .Z(n856) );
  IVSVTX2 U625 ( .A(n1883), .Z(n3773) );
  CTIVSVTX2 U626 ( .A(n3728), .Z(n585) );
  CTBUFSVTX2 U627 ( .A(n3215), .Z(n862) );
  CTIVSVTX4 U628 ( .A(n1422), .Z(n527) );
  IVSVTX0H U629 ( .A(n1790), .Z(n1315) );
  IVSVTX8 U630 ( .A(n1676), .Z(n3117) );
  NR2ASVTX6 U631 ( .A(n715), .B(n4023), .Z(n3622) );
  IVSVTX2 U632 ( .A(n1588), .Z(n1587) );
  ND2SVTX2 U633 ( .A(n4031), .B(n4030), .Z(n4041) );
  AN3SVTX2 U634 ( .A(n3712), .B(n3711), .C(n3710), .Z(n3713) );
  ND2SVTX2 U635 ( .A(n3155), .B(n3154), .Z(n1430) );
  ND2SVTX4 U636 ( .A(n3134), .B(n4159), .Z(n1279) );
  ND2SVTX2 U637 ( .A(n4066), .B(n487), .Z(n1103) );
  IVSVTX0H U638 ( .A(n3693), .Z(n3697) );
  ND2SVTX4 U639 ( .A(n1496), .B(n2010), .Z(n1495) );
  ND3SVTX2 U640 ( .A(n1386), .B(n3677), .C(n3676), .Z(n1385) );
  IVSVTX2 U641 ( .A(n1591), .Z(n1292) );
  AO7SVTX2 U642 ( .A(n3311), .B(n2378), .C(n4069), .Z(n3216) );
  IVSVTX1 U643 ( .A(n1474), .Z(n1657) );
  ND3SVTX4 U644 ( .A(n3884), .B(n446), .C(n3883), .Z(n2340) );
  IVSVTX2 U645 ( .A(n3333), .Z(n2025) );
  B_ND2SVTX2 U646 ( .A(n3897), .B(n3893), .Z(n2431) );
  NR2SVTX2 U647 ( .A(n3138), .B(n3139), .Z(n3141) );
  ND2SVTX4 U648 ( .A(n3917), .B(n3916), .Z(n3922) );
  F_ND3SVTX2 U649 ( .A(n3630), .B(n2067), .C(n3780), .Z(n2101) );
  ND4SVTX4 U650 ( .A(n1302), .B(n1303), .C(n1301), .D(n3178), .Z(n3185) );
  NR2SVTX2 U651 ( .A(n4163), .B(n4140), .Z(n4100) );
  OR2SVTX2 U652 ( .A(n4118), .B(n3202), .Z(n3210) );
  ND4SVTX4 U653 ( .A(n3739), .B(n1864), .C(n3634), .D(n3631), .Z(n3648) );
  ND2SVTX4 U654 ( .A(n486), .B(n4032), .Z(n2024) );
  F_IVSVTX1 U655 ( .A(n4139), .Z(n563) );
  AO6ASVTX2 U656 ( .A(n536), .B(n3998), .C(n1409), .Z(n3320) );
  AO7SVTX4 U657 ( .A(n3423), .B(n785), .C(n1488), .Z(n3426) );
  AO17ASVTX4 U658 ( .A(n1666), .B(n1314), .C(n1312), .D(n2292), .Z(n1311) );
  AO17SVTX6 U659 ( .A(n4022), .B(n3845), .C(n3844), .D(n3843), .Z(n1753) );
  B_ND2SVTX2 U660 ( .A(n3596), .B(n1690), .Z(n989) );
  NR3SVTX4 U661 ( .A(n2248), .B(n3184), .C(n3180), .Z(n3176) );
  CTIVSVTX2 U662 ( .A(n2424), .Z(n1293) );
  NR2ASVTX2 U663 ( .A(n593), .B(n3685), .Z(n1266) );
  ND2ASVTX4 U664 ( .A(n389), .B(n2103), .Z(n2071) );
  CTBUFSVTX8 U665 ( .A(n2352), .Z(n441) );
  NR2SVTX2 U666 ( .A(n3705), .B(n1824), .Z(n1428) );
  OR2SVTX2 U667 ( .A(n3247), .B(n3129), .Z(n3136) );
  NR2SVTX4 U668 ( .A(n526), .B(n1864), .Z(n3635) );
  NR3SVTX4 U669 ( .A(n587), .B(n3918), .C(n1740), .Z(n3919) );
  ND2ASVTX1 U670 ( .A(n3893), .B(n3898), .Z(n2080) );
  F_ENSVTX2 U671 ( .A(n506), .B(n2776), .Z(n4163) );
  IVSVTX6 U672 ( .A(n2360), .Z(n1697) );
  IVSVTX6 U673 ( .A(n961), .Z(n960) );
  IVSVTX6 U674 ( .A(n3742), .Z(n562) );
  ND2ASVTX6 U675 ( .A(n2929), .B(n1269), .Z(n1244) );
  IVSVTX0H U676 ( .A(n3880), .Z(n1666) );
  CTIVSVTX2 U677 ( .A(n3653), .Z(n515) );
  IVSVTX2 U678 ( .A(n1270), .Z(n3190) );
  IVSVTX2 U679 ( .A(n2140), .Z(n2139) );
  IVSVTX2 U680 ( .A(n3793), .Z(n3790) );
  BFSVTX10 U681 ( .A(n2393), .Z(n1705) );
  IVSVTX0H U682 ( .A(n3982), .Z(n753) );
  F_AN2SVTX2 U683 ( .A(n4014), .B(n2416), .Z(n3940) );
  IVSVTX0H U684 ( .A(n3372), .Z(n3373) );
  ND2SVTX4 U685 ( .A(n644), .B(n1499), .Z(n3903) );
  NR2ASVTX1 U686 ( .A(n593), .B(n3597), .Z(n3596) );
  CTIVSVTX2 U687 ( .A(n715), .Z(n1698) );
  IVSVTX4 U688 ( .A(n1329), .Z(n1328) );
  ND2SVTX2 U689 ( .A(n2801), .B(n780), .Z(n3351) );
  AN2SVTX4 U690 ( .A(n2442), .B(n3203), .Z(n3264) );
  IVSVTX2 U691 ( .A(n528), .Z(n1910) );
  NR2ASVTX4 U692 ( .A(n3871), .B(n3870), .Z(n3878) );
  IVSVTX4 U693 ( .A(n3613), .Z(n2248) );
  IVSVTX2 U694 ( .A(n1796), .Z(n2136) );
  ND2SVTX2 U695 ( .A(n1634), .B(n2352), .Z(n1140) );
  F_IVSVTX1 U696 ( .A(n3851), .Z(n3844) );
  B_ND2SVTX2 U697 ( .A(n3913), .B(n1658), .Z(n3917) );
  NR2SVTX4 U698 ( .A(n3977), .B(n3423), .Z(n3425) );
  BFSVTX8 U699 ( .A(n4171), .Z(n1596) );
  AO6ABSVTX4 U700 ( .A(n3332), .B(n3129), .C(n3128), .Z(n3134) );
  NR2ASVTX4 U701 ( .A(n530), .B(n3754), .Z(n3755) );
  ND2SVTX6 U702 ( .A(n3719), .B(n3795), .Z(n1417) );
  CTIVSVTX2 U703 ( .A(n3204), .Z(n3205) );
  ND2SVTX2 U704 ( .A(n770), .B(n3334), .Z(n1693) );
  NR2SVTX4 U705 ( .A(n2437), .B(n3371), .Z(n3333) );
  ND2ASVTX4 U706 ( .A(n534), .B(n486), .Z(n3251) );
  NR2SVTX2 U707 ( .A(n3609), .B(n1863), .Z(n3615) );
  AO7NSVTX4 U708 ( .A(n587), .B(n1740), .C(n3915), .Z(n3916) );
  ND2SVTX4 U709 ( .A(n705), .B(n1338), .Z(n3798) );
  ND3ABSVTX2 U710 ( .A(n3899), .B(n3898), .C(n679), .Z(n3900) );
  NR3ABSVTX4 U711 ( .A(n1864), .B(n533), .C(n3950), .Z(n3952) );
  ND2SVTX2 U712 ( .A(n1518), .B(n2103), .Z(n1196) );
  AO4SVTX4 U713 ( .A(n3666), .B(n2242), .C(n1824), .D(n2242), .Z(n1383) );
  AO1ABSVTX6 U714 ( .A(n3788), .B(n3740), .C(n526), .D(n3741), .Z(n1729) );
  ND4SVTX2 U715 ( .A(n3670), .B(n3672), .C(n3671), .D(n3669), .Z(n3677) );
  ND2SVTX4 U716 ( .A(n3114), .B(n4068), .Z(n1588) );
  ND2SVTX2 U717 ( .A(n4117), .B(n531), .Z(n1487) );
  NR2ASVTX2 U718 ( .A(n3912), .B(n2207), .Z(n2206) );
  F_ENSVTX2 U719 ( .A(n3556), .B(n3555), .Z(n3559) );
  FA1SVTX1 U720 ( .A(n3024), .B(n606), .CI(n3024), .Z(n2826) );
  ND2SVTX8 U721 ( .A(n1206), .B(n2914), .Z(n3893) );
  IVSVTX2 U722 ( .A(n3201), .Z(n4118) );
  IVSVTX6 U723 ( .A(n3686), .Z(n2067) );
  IVSVTX8 U724 ( .A(n991), .Z(n1635) );
  CTIVSVTX2 U725 ( .A(n3673), .Z(n1609) );
  IVSVTX2 U726 ( .A(n2393), .Z(n1854) );
  IVSVTX4 U727 ( .A(n3215), .Z(n2378) );
  CTIVSVTX2 U728 ( .A(n3710), .Z(n3666) );
  ND2SVTX4 U729 ( .A(n2938), .B(n2937), .Z(n1591) );
  ND2ASVTX4 U730 ( .A(n3122), .B(n3037), .Z(n3332) );
  IVSVTX0H U731 ( .A(n3603), .Z(n3639) );
  NR2ASVTX4 U732 ( .A(n3201), .B(n3206), .Z(n3150) );
  IVSVTX0H U733 ( .A(n3897), .Z(n3899) );
  IVSVTX8 U734 ( .A(n1863), .Z(n1864) );
  IVSVTX4 U735 ( .A(n4133), .Z(n3112) );
  IVSVTX2 U736 ( .A(n4158), .Z(n770) );
  B_ND2SVTX2 U737 ( .A(n3984), .B(n3983), .Z(n3987) );
  IVSVTX0H U738 ( .A(n4035), .Z(n3394) );
  ND2SVTX2 U739 ( .A(n3817), .B(n3681), .Z(n3633) );
  ND2SVTX6 U740 ( .A(n3928), .B(n2171), .Z(n1530) );
  IVSVTX2 U741 ( .A(n3973), .Z(n3423) );
  IVSVTX0H U742 ( .A(n3386), .Z(n3359) );
  IVSVTX2 U743 ( .A(n3929), .Z(n3950) );
  IVSVTX2 U744 ( .A(n3966), .Z(n1195) );
  IVSVTX2 U745 ( .A(n4010), .Z(n4012) );
  B_ND2SVTX2 U746 ( .A(n3656), .B(n3568), .Z(n3658) );
  F_IVSVTX1 U747 ( .A(n3914), .Z(n2207) );
  B_ND2SVTX2 U748 ( .A(n3783), .B(n2463), .Z(n3751) );
  AN2SVTX2 U749 ( .A(n3471), .B(n3557), .Z(n2464) );
  CTBUFSVTX6 U750 ( .A(n3855), .Z(n1658) );
  IVSVTX4 U751 ( .A(n765), .Z(n2103) );
  ND2ASVTX4 U752 ( .A(n697), .B(n475), .Z(n2247) );
  IVSVTX2 U753 ( .A(n3446), .Z(n3438) );
  F_ND2ASVTX2 U754 ( .A(n507), .B(n3396), .Z(n4031) );
  ENSVTX1 U755 ( .A(n3452), .B(n2746), .Z(n2380) );
  ND2SVTX2 U756 ( .A(n1993), .B(n2301), .Z(n3945) );
  MUX21NSVTX1 U757 ( .A(n3672), .B(n824), .S(n3671), .Z(n3674) );
  ENSVTX0H U758 ( .A(n3534), .B(n3535), .Z(n3536) );
  ND2SVTX4 U759 ( .A(n3787), .B(n3788), .Z(n3793) );
  ND2SVTX2 U760 ( .A(n3078), .B(n2352), .Z(n1213) );
  B_ND2SVTX2 U761 ( .A(n2296), .B(n535), .Z(n2422) );
  AO6CSVTX6 U762 ( .A(n388), .B(n2457), .C(n3911), .Z(n481) );
  IVSVTX4 U763 ( .A(n1473), .Z(n1474) );
  IVSVTX4 U764 ( .A(n4068), .Z(n1700) );
  AO7SVTX2 U765 ( .A(n2399), .B(n485), .C(n3882), .Z(n3881) );
  AO7SVTX4 U766 ( .A(n3464), .B(n405), .C(n1674), .Z(n404) );
  NR2SVTX2 U767 ( .A(n3544), .B(n3545), .Z(n1611) );
  BFSVTX2 U768 ( .A(n3981), .Z(n1885) );
  BFSVTX6 U769 ( .A(n3619), .Z(n880) );
  B_ND2SVTX2 U770 ( .A(n2416), .B(n4009), .Z(n1869) );
  ND3SVTX4 U771 ( .A(n4014), .B(n3939), .C(n3784), .Z(n3753) );
  ND2SVTX2 U772 ( .A(n3465), .B(n577), .Z(n1674) );
  CTBUFSVTX4 U773 ( .A(n3531), .Z(n373) );
  IVSVTX2 U774 ( .A(n3704), .Z(n1148) );
  ND2ASVTX6 U775 ( .A(n2941), .B(n2797), .Z(n3114) );
  OR2SVTX6 U776 ( .A(n2938), .B(n2937), .Z(n2393) );
  IVSVTX8 U777 ( .A(n1259), .Z(n1863) );
  F_ENSVTX2 U778 ( .A(n700), .B(n699), .Z(n698) );
  CTBUFSVTX4 U779 ( .A(n3391), .Z(n1321) );
  IVSVTX2 U780 ( .A(n3105), .Z(n1303) );
  IVSVTX2 U781 ( .A(n4121), .Z(n2949) );
  IVSVTX1 U782 ( .A(n2829), .Z(n3841) );
  CTIVSVTX2 U783 ( .A(n3872), .Z(n877) );
  CTIVSVTX2 U784 ( .A(n2050), .Z(n586) );
  F_AN2SVTX2 U785 ( .A(n3880), .B(n3865), .Z(n2399) );
  IVSVTX2 U786 ( .A(n1638), .Z(n3174) );
  B_ND2SVTX2 U787 ( .A(n3588), .B(n955), .Z(n3543) );
  NR2SVTX4 U788 ( .A(n3422), .B(n1079), .Z(n785) );
  B_ND2SVTX2 U789 ( .A(n3539), .B(n3589), .Z(n3545) );
  IVSVTX0H U790 ( .A(n3681), .Z(n3611) );
  ND2SVTX2 U791 ( .A(n1488), .B(n3973), .Z(n3974) );
  NR2SVTX6 U792 ( .A(n1354), .B(n1517), .Z(n1409) );
  ND3SVTX2 U793 ( .A(n3603), .B(n3641), .C(n3640), .Z(n3642) );
  ND2SVTX2 U794 ( .A(n3897), .B(n3764), .Z(n3856) );
  ND2ASVTX4 U795 ( .A(n510), .B(n3663), .Z(n3707) );
  IVSVTX2 U796 ( .A(n644), .Z(n1324) );
  IVSVTX2 U797 ( .A(n3680), .Z(n422) );
  ND3ASVTX4 U798 ( .A(n3084), .B(n3473), .C(n3472), .Z(n1218) );
  CTIVSVTX2 U799 ( .A(n3817), .Z(n3810) );
  AO6SVTX4 U800 ( .A(n4014), .B(n3889), .C(n3888), .Z(n3890) );
  AN2SVTX2 U801 ( .A(n492), .B(n3835), .Z(n3831) );
  ND2SVTX6 U802 ( .A(n3620), .B(n3619), .Z(n2065) );
  IVSVTX4 U803 ( .A(n3660), .Z(n1473) );
  NR2SVTX2 U804 ( .A(n3465), .B(n577), .Z(n3466) );
  AO7SVTX6 U805 ( .A(n1373), .B(n1122), .C(n3620), .Z(n3445) );
  IVSVTX0H U806 ( .A(n2347), .Z(n3281) );
  NR2SVTX2 U807 ( .A(n3463), .B(n3462), .Z(n3469) );
  IVSVTX2 U808 ( .A(n3795), .Z(n3797) );
  AN2SVTX4 U809 ( .A(n2416), .B(n1991), .Z(n1994) );
  IVSVTX4 U810 ( .A(n3920), .Z(n388) );
  NR2ASVTX6 U811 ( .A(n3764), .B(n3413), .Z(n3983) );
  IVSVTX2 U812 ( .A(n2920), .Z(n2913) );
  ND2SVTX4 U813 ( .A(n3764), .B(n3885), .Z(n3898) );
  IVSVTX2 U814 ( .A(n3927), .Z(n4001) );
  CTIVSVTX2 U815 ( .A(n2825), .Z(n1354) );
  ND2ASVTX6 U816 ( .A(n505), .B(n3661), .Z(n3710) );
  IVSVTX2 U817 ( .A(n3484), .Z(n3485) );
  IVSVTX10 U818 ( .A(n2292), .Z(n3686) );
  EN3SVTX6 U819 ( .A(n342), .B(n1571), .C(n622), .Z(n1923) );
  IVSVTX2 U820 ( .A(n1299), .Z(n3874) );
  NR2ASVTX4 U821 ( .A(n516), .B(n3310), .Z(n930) );
  IVSVTX2 U822 ( .A(n3930), .Z(n3931) );
  IVSVTX2 U823 ( .A(n2935), .Z(n2163) );
  CTBUFSVTX4 U824 ( .A(n3933), .Z(n415) );
  IVSVTX2 U825 ( .A(n2946), .Z(n2290) );
  IVSVTX2 U826 ( .A(n3472), .Z(n3476) );
  CTIVSVTX4 U827 ( .A(n3621), .Z(n511) );
  ND2SVTX2 U828 ( .A(n3816), .B(n3817), .Z(n2452) );
  NR2ASVTX4 U829 ( .A(n3544), .B(n3538), .Z(n3498) );
  ND2SVTX2 U830 ( .A(n2987), .B(n2763), .Z(n700) );
  ENSVTX1 U831 ( .A(n3518), .B(n3517), .Z(n702) );
  ND2SVTX2 U832 ( .A(n2327), .B(n3025), .Z(n3028) );
  B_ND2SVTX2 U833 ( .A(n2866), .B(n2867), .Z(n3165) );
  NR2SVTX2 U834 ( .A(n601), .B(n1655), .Z(n346) );
  ND2SVTX2 U835 ( .A(n3471), .B(n3458), .Z(n3463) );
  CTIVSVTX2 U836 ( .A(n3764), .Z(n3414) );
  ND2SVTX4 U837 ( .A(n3571), .B(n3572), .Z(n1066) );
  IVSVTX2 U838 ( .A(n742), .Z(n1364) );
  ND2ASVTX4 U839 ( .A(n510), .B(n1146), .Z(n1511) );
  NR2SVTX6 U840 ( .A(n2920), .B(n3981), .Z(n1203) );
  ND2ASVTX4 U841 ( .A(n389), .B(n1902), .Z(n3926) );
  NR3SVTX6 U842 ( .A(n3048), .B(n1319), .C(n3105), .Z(n1982) );
  B_ND2SVTX2 U843 ( .A(n2933), .B(n2934), .Z(n2162) );
  CTIVSVTX2 U844 ( .A(n833), .Z(n2824) );
  ND2SVTX2 U845 ( .A(n3097), .B(n3096), .Z(n3737) );
  IVSVTX2 U846 ( .A(n609), .Z(n2385) );
  CTIVSVTX2 U847 ( .A(n2773), .Z(n2774) );
  ND2ASVTX6 U848 ( .A(n3570), .B(n3443), .Z(n3571) );
  BFSVTX4 U849 ( .A(n1327), .Z(n3684) );
  IVSVTX2 U850 ( .A(n610), .Z(n516) );
  IVSVTX2 U851 ( .A(n2921), .Z(n2873) );
  CTIVSVTX2 U852 ( .A(n3980), .Z(n590) );
  IVSVTX2 U853 ( .A(n713), .Z(n1856) );
  B_ND2SVTX2 U854 ( .A(n1766), .B(n3483), .Z(n2244) );
  IVSVTX4 U855 ( .A(n2198), .Z(n2200) );
  IVSVTX2 U856 ( .A(n2379), .Z(n584) );
  CTAN2BSVTX4 U857 ( .A(n1518), .B(n623), .Z(n3749) );
  CTIVSVTX2 U858 ( .A(n3607), .Z(n3608) );
  IVSVTX4 U859 ( .A(n2077), .Z(n2457) );
  NR2ASVTX2 U860 ( .A(n1518), .B(n539), .Z(n3935) );
  IVSVTX4 U861 ( .A(n3912), .Z(n587) );
  ND2SVTX6 U862 ( .A(n2179), .B(n833), .Z(n1902) );
  IVSVTX0H U863 ( .A(n3887), .Z(n755) );
  IVSVTX2 U864 ( .A(n3411), .Z(n2912) );
  AO7SVTX4 U865 ( .A(n3526), .B(n2420), .C(n3525), .Z(n3572) );
  CTIVSVTX2 U866 ( .A(n955), .Z(n3538) );
  NR2SVTX2 U867 ( .A(n3091), .B(n3088), .Z(n3092) );
  IVSVTX2 U868 ( .A(n3818), .Z(n3811) );
  NR2SVTX2 U869 ( .A(n3096), .B(n3097), .Z(n3052) );
  IVSVTX4 U870 ( .A(n1271), .Z(n742) );
  ND2SVTX4 U871 ( .A(n2909), .B(n2908), .Z(n3911) );
  ND2SVTX2 U872 ( .A(n3963), .B(n485), .Z(n1830) );
  F_ENSVTX2 U873 ( .A(n1788), .B(n3122), .Z(n3008) );
  CTIVSVTX2 U874 ( .A(n2339), .Z(n1366) );
  NR2ASVTX2 U875 ( .A(n2971), .B(n1347), .Z(n3746) );
  ND2ASVTX6 U876 ( .A(n3061), .B(n3088), .Z(n3809) );
  ND2ASVTX6 U877 ( .A(n517), .B(n3449), .Z(n3519) );
  ND2ASVTX6 U878 ( .A(n2821), .B(n1019), .Z(n3840) );
  CTIVSVTX6 U879 ( .A(n3122), .Z(n507) );
  EO3SVTX6 U880 ( .A(n3311), .B(n1334), .C(n2185), .Z(n1517) );
  IVSVTX2 U881 ( .A(n3586), .Z(n2325) );
  ND2SVTX4 U882 ( .A(n2916), .B(n2915), .Z(n3885) );
  ND2ASVTX6 U883 ( .A(n607), .B(n2877), .Z(n3702) );
  ND2SVTX4 U884 ( .A(n2880), .B(n2881), .Z(n3704) );
  NR2ASVTX4 U885 ( .A(n1149), .B(n2883), .Z(n3451) );
  B_ND2SVTX2 U886 ( .A(n1030), .B(n1881), .Z(n3667) );
  NR2ASVTX2 U887 ( .A(n503), .B(n624), .Z(n2462) );
  B_ND2SVTX2 U888 ( .A(n2925), .B(n2924), .Z(n3224) );
  ND2SVTX6 U889 ( .A(n3566), .B(n2372), .Z(n3568) );
  ENSVTX6 U890 ( .A(n3038), .B(n1242), .Z(n3310) );
  F_ND2ASVTX2 U891 ( .A(n2971), .B(n1347), .Z(n3748) );
  ND2SVTX6 U892 ( .A(n3607), .B(n3606), .Z(n3808) );
  IVSVTX2 U893 ( .A(n1963), .Z(n1962) );
  CTIVSVTX4 U894 ( .A(n1835), .Z(n1344) );
  ND2SVTX6 U895 ( .A(n1450), .B(n2845), .Z(n2066) );
  IVSVTX2 U896 ( .A(n3483), .Z(n1633) );
  ND2SVTX6 U897 ( .A(n1204), .B(n2339), .Z(n3411) );
  CTIVSVTX2 U898 ( .A(n3102), .Z(n3103) );
  F_ENSVTX2 U899 ( .A(n506), .B(n2868), .Z(n2928) );
  AO5SVTX4 U900 ( .A(n1547), .B(n1932), .C(n624), .Z(n3022) );
  ND2ASVTX4 U901 ( .A(n1786), .B(n3584), .Z(n3963) );
  NR2SVTX2 U902 ( .A(n602), .B(n3886), .Z(n1870) );
  AO7SVTX6 U903 ( .A(n3552), .B(n1261), .C(n3550), .Z(n1823) );
  AO6SVTX2 U904 ( .A(n3042), .B(n3044), .C(n3043), .Z(n3045) );
  AN2SVTX4 U905 ( .A(n1730), .B(n539), .Z(n4007) );
  CTIVSVTX2 U906 ( .A(n2818), .Z(n1342) );
  ND2SVTX2 U907 ( .A(n2807), .B(n3122), .Z(n1793) );
  CTBUFSVTX4 U908 ( .A(n2017), .Z(n402) );
  IVSVTX2 U909 ( .A(n3005), .Z(n2965) );
  IVSVTX2 U910 ( .A(n1551), .Z(n727) );
  ND2ASVTX6 U911 ( .A(n517), .B(n3433), .Z(n3518) );
  IVSVTX2 U912 ( .A(n3503), .Z(n1606) );
  IVSVTX4 U913 ( .A(n2799), .Z(n2800) );
  CTIVSVTX2 U914 ( .A(n2876), .Z(n2877) );
  EN3SVTX6 U915 ( .A(n2788), .B(n948), .C(n621), .Z(n2961) );
  ND2ASVTX6 U916 ( .A(n1717), .B(n1634), .Z(n3532) );
  IVSVTX6 U917 ( .A(n1024), .Z(n1766) );
  IVSVTX2 U918 ( .A(n2719), .Z(n2726) );
  ND2SVTX2 U919 ( .A(n3626), .B(n3583), .Z(n1594) );
  B_ND2SVTX2 U920 ( .A(n3283), .B(n1030), .Z(n3478) );
  NR2ASVTX2 U921 ( .A(n2784), .B(n2945), .Z(n1257) );
  ND2SVTX4 U922 ( .A(n2419), .B(n3551), .Z(n3550) );
  IVSVTX4 U923 ( .A(n2845), .Z(n1436) );
  B_ND2SVTX2 U924 ( .A(n3494), .B(n3516), .Z(n3435) );
  IVSVTX2 U925 ( .A(n2879), .Z(n1062) );
  IVSVTX2 U926 ( .A(n1978), .Z(n1206) );
  AN2SVTX2 U927 ( .A(n814), .B(n2971), .Z(n3828) );
  ND2SVTX4 U928 ( .A(n2874), .B(n2875), .Z(n2925) );
  AN2SVTX2 U929 ( .A(n546), .B(n2858), .Z(n484) );
  ND3ASVTX6 U930 ( .A(n802), .B(n3460), .C(n3458), .Z(n804) );
  CTIVSVTX2 U931 ( .A(n1518), .Z(n1730) );
  CTIVSVTX4 U932 ( .A(n3625), .Z(n1711) );
  CTIVSVTX4 U933 ( .A(n1169), .Z(n1171) );
  B_ND2SVTX2 U934 ( .A(n2149), .B(n1695), .Z(n2347) );
  AN2SVTX4 U935 ( .A(n2815), .B(n2816), .Z(n1800) );
  ND2SVTX2 U936 ( .A(n2871), .B(n2870), .Z(n2922) );
  NR4SVTX6 U937 ( .A(n2776), .B(n2297), .C(n2722), .D(n2723), .Z(n1867) );
  ND2SVTX2 U938 ( .A(n390), .B(n1526), .Z(n1333) );
  AO7CSVTX2 U939 ( .A(n2807), .B(n3122), .C(n1006), .Z(n1792) );
  ND2ASVTX4 U940 ( .A(n1964), .B(n824), .Z(n1963) );
  ND3SVTX4 U941 ( .A(n3818), .B(n3816), .C(n3817), .Z(n3064) );
  AO5SVTX4 U942 ( .A(n1655), .B(n601), .C(n3880), .Z(n2020) );
  IVSVTX2 U943 ( .A(n623), .Z(n2223) );
  CTBUFSVTX4 U944 ( .A(n948), .Z(n444) );
  CTIVSVTX2 U945 ( .A(n2816), .Z(n1691) );
  EO3SVTX6 U946 ( .A(n3271), .B(n1361), .C(n1791), .Z(n2908) );
  IVSVTX2 U947 ( .A(n2923), .Z(n1168) );
  BFSVTX0H U948 ( .A(n1121), .Z(n1695) );
  EOSVTX1 U949 ( .A(n3279), .B(n3065), .Z(n456) );
  CTIVSVTX2 U950 ( .A(n2893), .Z(n2879) );
  IVSVTX2 U951 ( .A(n2815), .Z(n1692) );
  IVSVTX2 U952 ( .A(n2980), .Z(n2189) );
  IVSVTX4 U953 ( .A(n3723), .Z(n600) );
  ND2SVTX2 U954 ( .A(n3067), .B(n3283), .Z(n3493) );
  ND2ASVTX4 U955 ( .A(n1939), .B(n508), .Z(n3516) );
  ND2SVTX2 U956 ( .A(n2776), .B(n3024), .Z(n2727) );
  ND2ASVTX6 U957 ( .A(n2887), .B(n2762), .Z(n2763) );
  BFSVTX8 U958 ( .A(n1759), .Z(n1571) );
  AO7SVTX2 U959 ( .A(n2971), .B(n3311), .C(n1347), .Z(n1681) );
  ND2SVTX2 U960 ( .A(n823), .B(n1397), .Z(n3603) );
  ND2SVTX6 U961 ( .A(n841), .B(n840), .Z(n1551) );
  IVSVTX4 U962 ( .A(n3456), .Z(n1943) );
  ND2SVTX6 U963 ( .A(n3001), .B(n3000), .Z(n3489) );
  B_ND2SVTX2 U964 ( .A(n1892), .B(n1330), .Z(n1332) );
  OR2BSVTX4 U965 ( .A(n537), .B(n3068), .Z(n3636) );
  ND2SVTX2 U966 ( .A(n3827), .B(n3887), .Z(n3289) );
  ND2SVTX2 U967 ( .A(n2149), .B(n2843), .Z(n2169) );
  IVSVTX6 U968 ( .A(n540), .Z(n2868) );
  ND3SVTX4 U969 ( .A(n616), .B(n2720), .C(n3126), .Z(n2723) );
  IVSVTX4 U970 ( .A(n3471), .Z(n3084) );
  ND2SVTX2 U971 ( .A(n3122), .B(n3311), .Z(n2874) );
  IVSVTX2 U972 ( .A(n2387), .Z(n1983) );
  NR2ASVTX1 U973 ( .A(n543), .B(n969), .Z(n2852) );
  AO7SVTX6 U974 ( .A(n1932), .B(n615), .C(n432), .Z(n1232) );
  NR2SVTX6 U975 ( .A(n2419), .B(n3551), .Z(n1261) );
  AO7SVTX6 U976 ( .A(n3043), .B(n3042), .C(n3044), .Z(n1320) );
  F_ENSVTX2 U977 ( .A(n1268), .B(n3079), .Z(n1828) );
  ENSVTX4 U978 ( .A(n621), .B(n779), .Z(n1169) );
  AN2SVTX2 U979 ( .A(n623), .B(n396), .Z(n3051) );
  IVSVTX8 U980 ( .A(n1295), .Z(n1932) );
  IVSVTX6 U981 ( .A(n3126), .Z(n3111) );
  IVSVTX2 U982 ( .A(n997), .Z(n996) );
  EO3SVTX6 U983 ( .A(n3065), .B(n1647), .C(n1851), .Z(n2892) );
  ND2ASVTX4 U984 ( .A(n2814), .B(n2168), .Z(n2191) );
  AO7CSVTX4 U985 ( .A(n2905), .B(n728), .C(n1347), .Z(n398) );
  CTBUFSVTX4 U986 ( .A(n1346), .Z(n342) );
  IVSVTX2 U987 ( .A(n1764), .Z(n396) );
  IVSVTX10 U988 ( .A(n2788), .Z(n615) );
  CTIVSVTX6 U989 ( .A(n3000), .Z(n1758) );
  ND2ASVTX6 U990 ( .A(n911), .B(n686), .Z(n3494) );
  IVSVTX10 U991 ( .A(n3126), .Z(n3122) );
  IVSVTX4 U992 ( .A(n539), .Z(n1789) );
  CTBUFSVTX4 U993 ( .A(n518), .Z(n432) );
  ND2ASVTX6 U994 ( .A(n473), .B(n1709), .Z(n3001) );
  IVSVTX2 U995 ( .A(n2973), .Z(n2975) );
  IVSVTX4 U996 ( .A(n2807), .Z(n1728) );
  IVSVTX6 U997 ( .A(n3958), .Z(n1335) );
  IVSVTX6 U998 ( .A(n2789), .Z(n606) );
  ND2SVTX2 U999 ( .A(n1223), .B(n1791), .Z(n2906) );
  ND2SVTX4 U1000 ( .A(n1547), .B(n622), .Z(n760) );
  IVSVTX2 U1001 ( .A(n728), .Z(n520) );
  IVSVTX4 U1002 ( .A(n2822), .Z(n1664) );
  B_ND2SVTX2 U1003 ( .A(n612), .B(n997), .Z(n995) );
  IVSVTX4 U1004 ( .A(n2974), .Z(n2300) );
  ND2ASVTX4 U1005 ( .A(n684), .B(n538), .Z(n3285) );
  F_ND2ASVTX2 U1006 ( .A(n2998), .B(n2999), .Z(n1809) );
  AO7SVTX4 U1007 ( .A(n1482), .B(n1518), .C(n948), .Z(n772) );
  BFSVTX1 U1008 ( .A(n1937), .Z(n1601) );
  AO17ASVTX4 U1009 ( .A(n630), .B(n508), .C(n687), .D(n3286), .Z(n2882) );
  AO5SVTX2 U1010 ( .A(n1295), .B(n503), .C(n2971), .Z(n2897) );
  F_ND2ASVTX1 U1011 ( .A(n630), .B(n3065), .Z(n1150) );
  F_ND2ASVTX2 U1012 ( .A(n2398), .B(n1518), .Z(n2037) );
  F_ENSVTX2 U1013 ( .A(n1717), .B(n684), .Z(n2762) );
  F_ND2ASVTX2 U1014 ( .A(n1881), .B(n2814), .Z(n3638) );
  IVSVTX6 U1015 ( .A(n357), .Z(n2835) );
  BFSVTX12 U1016 ( .A(n4018), .Z(n1347) );
  CTBUFSVTX4 U1017 ( .A(n617), .Z(n390) );
  IVSVTX6 U1018 ( .A(n2398), .Z(n1482) );
  BFSVTX6 U1019 ( .A(n3065), .Z(n428) );
  BFSVTX8 U1020 ( .A(n625), .Z(n1686) );
  IVSVTX2 U1021 ( .A(n2888), .Z(n2885) );
  IVSVTX2 U1022 ( .A(n3279), .Z(n969) );
  IVSVTX6 U1023 ( .A(n2348), .Z(n610) );
  IVSVTX2 U1024 ( .A(n2820), .Z(n2813) );
  BFSVTX8 U1025 ( .A(n2398), .Z(n624) );
  AO7SVTX2 U1026 ( .A(n1361), .B(n1339), .C(n3068), .Z(n2130) );
  BFSVTX4 U1027 ( .A(n2375), .Z(n2092) );
  ND2SVTX2 U1028 ( .A(n1361), .B(n502), .Z(n2978) );
  ND2SVTX2 U1029 ( .A(n608), .B(n3270), .Z(n2967) );
  IVSVTX6 U1030 ( .A(n2990), .Z(n2283) );
  BFSVTX8 U1031 ( .A(n3271), .Z(n1743) );
  ND2ASVTX4 U1032 ( .A(n2760), .B(n3079), .Z(n3286) );
  IVSVTX4 U1033 ( .A(n1251), .Z(n1254) );
  ND2SVTX6 U1034 ( .A(n2944), .B(n3024), .Z(n2743) );
  IVSVTX4 U1035 ( .A(n2995), .Z(n2992) );
  AO5SVTX4 U1036 ( .A(n1881), .B(n2151), .C(n625), .Z(n3091) );
  AO6SVTX4 U1037 ( .A(n2112), .B(n547), .C(n730), .Z(n1472) );
  AO7SVTX6 U1038 ( .A(n1006), .B(n539), .C(n617), .Z(n1355) );
  ND2SVTX4 U1039 ( .A(n2971), .B(n823), .Z(n1208) );
  AO7SVTX4 U1040 ( .A(n964), .B(n1481), .C(n1669), .Z(n1709) );
  ND3SVTX4 U1041 ( .A(n1030), .B(n3065), .C(n1669), .Z(n2733) );
  IVSVTX4 U1042 ( .A(n1529), .Z(n1143) );
  ND2SVTX2 U1043 ( .A(n1748), .B(n2032), .Z(n1049) );
  ENSVTX4 U1044 ( .A(n659), .B(n686), .Z(n2883) );
  ND2ASVTX4 U1045 ( .A(n3065), .B(n1618), .Z(n1151) );
  BFSVTX4 U1046 ( .A(n1939), .Z(n1634) );
  ND2ASVTX6 U1047 ( .A(n3032), .B(n2344), .Z(n2717) );
  IVSVTX2 U1048 ( .A(n541), .Z(n1741) );
  IVSVTX8 U1049 ( .A(n542), .Z(n2348) );
  ND2SVTX2 U1050 ( .A(n2784), .B(n2255), .Z(n2722) );
  IVSVTX2 U1051 ( .A(n2147), .Z(n919) );
  ND2SVTX2 U1052 ( .A(n1361), .B(n539), .Z(n1363) );
  B_ND2SVTX2 U1053 ( .A(n543), .B(n684), .Z(n2989) );
  AN2SVTX4 U1054 ( .A(n546), .B(n808), .Z(n2970) );
  F_ND2ASVTX2 U1055 ( .A(n2760), .B(n3065), .Z(n3074) );
  F_ENSVTX2 U1056 ( .A(n1480), .B(n626), .Z(n2150) );
  ND2SVTX4 U1057 ( .A(n2017), .B(n537), .Z(n1837) );
  BFSVTX4 U1058 ( .A(n3279), .Z(n1972) );
  IVSVTX4 U1059 ( .A(n391), .Z(n2731) );
  BFSVTX8 U1060 ( .A(n1529), .Z(n1526) );
  IVSVTX2 U1061 ( .A(n1748), .Z(n399) );
  IVSVTX2 U1062 ( .A(n1939), .Z(n1523) );
  BFSVTX10 U1063 ( .A(n2812), .Z(n942) );
  IVSVTX10 U1064 ( .A(n3273), .Z(n948) );
  CTIVSVTX6 U1065 ( .A(n3067), .Z(n538) );
  BFSVTX8 U1066 ( .A(n1199), .Z(n728) );
  CTBUFSVTX6 U1067 ( .A(n1121), .Z(n1618) );
  ND2SVTX2 U1068 ( .A(n2899), .B(n418), .Z(n2900) );
  F_ND2ASVTX2 U1069 ( .A(n543), .B(n546), .Z(n1827) );
  IVSVTX4 U1070 ( .A(n1748), .Z(n2151) );
  IVSVTX4 U1071 ( .A(n1529), .Z(n359) );
  IVSVTX6 U1072 ( .A(n1268), .Z(n543) );
  BFSVTX6 U1073 ( .A(n1025), .Z(n1042) );
  ND2ASVTX6 U1074 ( .A(n709), .B(n2240), .Z(n2284) );
  IVSVTX8 U1075 ( .A(n798), .Z(n3282) );
  BFSVTX6 U1076 ( .A(n1267), .Z(n1973) );
  IVSVTX10 U1077 ( .A(n500), .Z(n501) );
  F_ND2ASVTX2 U1078 ( .A(n1861), .B(n2751), .Z(n1860) );
  IVSVTX6 U1079 ( .A(n2282), .Z(n1701) );
  IVSVTX10 U1080 ( .A(n544), .Z(n709) );
  IVSVTX6 U1081 ( .A(n1358), .Z(n1480) );
  ND3SVTX6 U1082 ( .A(n2619), .B(n1287), .C(n2415), .Z(n1272) );
  B_ND2SVTX2 U1083 ( .A(n2601), .B(n2602), .Z(n1273) );
  ND3SVTX4 U1084 ( .A(n2600), .B(n776), .C(n820), .Z(n1274) );
  MUX21NSVTX6 U1085 ( .A(n2599), .B(n2269), .S(n631), .Z(n2899) );
  CTBUFSVTX4 U1086 ( .A(n2331), .Z(n338) );
  IVSVTX2 U1087 ( .A(n1124), .Z(n918) );
  IVSVTX10 U1088 ( .A(n798), .Z(n544) );
  IVSVTX6 U1089 ( .A(n1152), .Z(n1154) );
  IVSVTX8 U1090 ( .A(n683), .Z(n684) );
  IVSVTX2 U1091 ( .A(n2676), .Z(n1651) );
  IVSVTX4 U1092 ( .A(n915), .Z(n1965) );
  ND3SVTX6 U1093 ( .A(n2600), .B(n1287), .C(n1114), .Z(n786) );
  ND3SVTX6 U1094 ( .A(n2601), .B(n2602), .C(n776), .Z(n2596) );
  B_ND2SVTX2 U1095 ( .A(n2691), .B(n2692), .Z(n1605) );
  AO2ASVTX6 U1096 ( .C(n1043), .D(n2627), .A(n2668), .B(n2678), .Z(n675) );
  AO7SVTX6 U1097 ( .A(n2559), .B(n2558), .C(n2751), .Z(n1895) );
  CTBUFSVTX4 U1098 ( .A(n549), .Z(n418) );
  F_IVSVTX1 U1099 ( .A(n2593), .Z(n2548) );
  ND2SVTX4 U1100 ( .A(n1166), .B(n2982), .Z(n1165) );
  NR3SVTX4 U1101 ( .A(n2270), .B(n1287), .C(n2269), .Z(n1001) );
  ND3SVTX6 U1102 ( .A(n2655), .B(n2678), .C(n1210), .Z(n915) );
  ND2SVTX6 U1103 ( .A(n2839), .B(n632), .Z(n1886) );
  NR2SVTX2 U1104 ( .A(n2653), .B(n2652), .Z(n1893) );
  ND4SVTX4 U1105 ( .A(n707), .B(n2549), .C(n2550), .D(n680), .Z(n998) );
  ND2SVTX6 U1106 ( .A(n2587), .B(n1039), .Z(n776) );
  ND2SVTX2 U1107 ( .A(n891), .B(n2672), .Z(n2600) );
  BFSVTX8 U1108 ( .A(n1872), .Z(n1656) );
  ND2ASVTX6 U1109 ( .A(n2898), .B(n1039), .Z(n2616) );
  CTIVSVTX6 U1110 ( .A(n1026), .Z(n680) );
  CTBUFSVTX4 U1111 ( .A(n2618), .Z(n650) );
  IVSVTX2 U1112 ( .A(n549), .Z(n2270) );
  IVSVTX4 U1113 ( .A(n2110), .Z(n2599) );
  IVSVTX4 U1114 ( .A(n2654), .Z(n2269) );
  ND3ABSVTX4 U1115 ( .A(n2478), .B(n1107), .C(n1360), .Z(n2605) );
  IVSVTX4 U1116 ( .A(n2543), .Z(n2559) );
  IVSVTX4 U1117 ( .A(n1178), .Z(n2322) );
  ND2SVTX6 U1118 ( .A(n1287), .B(n2667), .Z(n692) );
  IVSVTX4 U1119 ( .A(n1116), .Z(n1894) );
  ND2ASVTX4 U1120 ( .A(n2668), .B(n2279), .Z(n685) );
  ND2SVTX4 U1121 ( .A(n2587), .B(n2610), .Z(n2591) );
  AO6SVTX4 U1122 ( .A(n2678), .B(n2671), .C(n2673), .Z(n2675) );
  ND2ASVTX6 U1123 ( .A(n1124), .B(n1127), .Z(n1119) );
  ND2SVTX4 U1124 ( .A(n2238), .B(n1060), .Z(n1167) );
  ND3SVTX6 U1125 ( .A(n2636), .B(n1233), .C(n1297), .Z(n1210) );
  IVSVTX2 U1126 ( .A(n2672), .Z(n2673) );
  ND2SVTX4 U1127 ( .A(n2700), .B(n2587), .Z(n682) );
  CTIVSVTX2 U1128 ( .A(n1116), .Z(n341) );
  NR2ASVTX2 U1129 ( .A(n2698), .B(n2697), .Z(n2699) );
  ND2ASVTX4 U1130 ( .A(n1107), .B(n2110), .Z(n2543) );
  CTIVSVTX2 U1131 ( .A(n2580), .Z(n416) );
  CTIVSVTX8 U1132 ( .A(n1115), .Z(n2279) );
  NR2SVTX2 U1133 ( .A(n550), .B(n1219), .Z(n653) );
  AO7SVTX2 U1134 ( .A(n2666), .B(n1360), .C(n2665), .Z(n2667) );
  AO7ASVTX4 U1135 ( .A(n2513), .B(n374), .C(n378), .Z(n655) );
  IVSVTX4 U1136 ( .A(n1872), .Z(n738) );
  IVSVTX10 U1137 ( .A(n1124), .Z(n1166) );
  BFSVTX0H U1138 ( .A(n2486), .Z(n378) );
  IVSVTX2 U1139 ( .A(n2563), .Z(n2314) );
  IVSVTX2 U1140 ( .A(n2184), .Z(n665) );
  CTBUFSVTX4 U1141 ( .A(n2652), .Z(n403) );
  BFSVTX0H U1142 ( .A(n2133), .Z(n2132) );
  IVSVTX4 U1143 ( .A(n1360), .Z(n968) );
  ND3SVTX6 U1144 ( .A(n1769), .B(n2579), .C(n2232), .Z(n2536) );
  CTBUFSVTX2 U1145 ( .A(n2503), .Z(n374) );
  NR2SVTX2 U1146 ( .A(n2589), .B(n2126), .Z(n1095) );
  ND2SVTX4 U1147 ( .A(n2566), .B(n2567), .Z(n693) );
  CTBUFSVTX4 U1148 ( .A(n2651), .Z(n857) );
  AO7SVTX1 U1149 ( .A(n2621), .B(n2574), .C(n639), .Z(n2081) );
  IVSVTX4 U1150 ( .A(n2618), .Z(n2036) );
  ND2ASVTX6 U1151 ( .A(n1117), .B(n512), .Z(n2898) );
  IVSVTX2 U1152 ( .A(n2651), .Z(n2323) );
  BFSVTX0H U1153 ( .A(n2577), .Z(n1629) );
  IVSVTX1 U1154 ( .A(n2671), .Z(n552) );
  ND2SVTX6 U1155 ( .A(n1112), .B(n1061), .Z(n2618) );
  ND2SVTX4 U1156 ( .A(n2638), .B(n1756), .Z(n2629) );
  IVSVTX0H U1157 ( .A(n920), .Z(n1861) );
  CTBUFSVTX2 U1158 ( .A(n963), .Z(n2572) );
  ND2ASVTX4 U1159 ( .A(n1723), .B(n2245), .Z(n2606) );
  F_ND2ASVTX2 U1160 ( .A(n553), .B(n513), .Z(n2312) );
  NR2ASVTX2 U1161 ( .A(n1035), .B(n1768), .Z(n1036) );
  IVSVTX10 U1162 ( .A(n1061), .Z(n1872) );
  IVSVTX2 U1163 ( .A(n2659), .Z(n2660) );
  BFSVTX6 U1164 ( .A(n2634), .Z(n2180) );
  IVSVTX0H U1165 ( .A(n551), .Z(n1035) );
  AN2SVTX4 U1166 ( .A(n2644), .B(n513), .Z(n2395) );
  IVSVTX10 U1167 ( .A(n1061), .Z(n1359) );
  IVSVTX2 U1168 ( .A(n2585), .Z(n431) );
  ND3SVTX6 U1169 ( .A(n2624), .B(n2232), .C(n1769), .Z(n1610) );
  ND2ASVTX4 U1170 ( .A(n2631), .B(n2561), .Z(n1767) );
  ND2SVTX2 U1171 ( .A(n2698), .B(n513), .Z(n846) );
  CTIVSVTX2 U1172 ( .A(n1545), .Z(n410) );
  IVSVTX2 U1173 ( .A(n2545), .Z(n2391) );
  IVSVTX2 U1174 ( .A(n2638), .Z(n635) );
  IVSVTX2 U1175 ( .A(num_i[3]), .Z(n555) );
  BFSVTX2 U1176 ( .A(num_i[9]), .Z(n2644) );
  IVSVTX10 U1177 ( .A(n2126), .Z(n1544) );
  IVSVTX10 U1178 ( .A(n2582), .Z(n1197) );
  IVSVTX2 U1179 ( .A(n2515), .Z(n1126) );
  IVSVTX2 U1180 ( .A(n393), .Z(n2512) );
  ND2SVTX4 U1181 ( .A(n1675), .B(n2544), .Z(n1936) );
  AN3SVTX4 U1182 ( .A(n2513), .B(n551), .C(n2377), .Z(n460) );
  IVSVTX4 U1183 ( .A(n2620), .Z(n2621) );
  NR2SVTX2 U1184 ( .A(n2588), .B(n2468), .Z(n1806) );
  IVSVTX4 U1185 ( .A(n1755), .Z(n551) );
  NR3SVTX4 U1186 ( .A(n2696), .B(n2695), .C(n2534), .Z(n2467) );
  IVSVTX6 U1187 ( .A(n2526), .Z(n2509) );
  IVSVTX4 U1188 ( .A(n658), .Z(n672) );
  CTBUFSVTX4 U1189 ( .A(num_i[23]), .Z(n891) );
  IVSVTX2 U1190 ( .A(num_i[9]), .Z(n2527) );
  BFSVTX2 U1191 ( .A(num_i[16]), .Z(n2588) );
  F_IVSVTX1 U1192 ( .A(n2518), .Z(n2369) );
  ND2SVTX6 U1193 ( .A(n1198), .B(n2499), .Z(n658) );
  ND3ASVTX6 U1194 ( .A(num_i[27]), .B(n2493), .C(n636), .Z(n2496) );
  IVSVTX8 U1195 ( .A(n2584), .Z(n636) );
  IVSVTX6 U1196 ( .A(n2534), .Z(n2578) );
  CTBUFSVTX4 U1197 ( .A(num_i[21]), .Z(n2696) );
  BFSVTX6 U1198 ( .A(num_i[19]), .Z(n2573) );
  NR2SVTX4 U1199 ( .A(num_i[16]), .B(num_i[19]), .Z(n2493) );
  NR2SVTX4 U1200 ( .A(num_i[27]), .B(num_i[28]), .Z(n1479) );
  NR2SVTX4 U1201 ( .A(num_i[18]), .B(num_i[16]), .Z(n2474) );
  NR2SVTX4 U1202 ( .A(num_i[30]), .B(num_i[29]), .Z(n2473) );
  IVSVTX8 U1203 ( .A(num_i[28]), .Z(n2577) );
  NR2SVTX6 U1204 ( .A(num_i[14]), .B(num_i[13]), .Z(n1031) );
  IVSVTX4 U1205 ( .A(n1209), .Z(n2228) );
  IVSVTX8 U1206 ( .A(n1085), .Z(n3443) );
  AO7ABSVTX2 U1207 ( .A(n543), .B(n508), .C(n2844), .Z(n714) );
  ND2SVTX2 U1208 ( .A(n628), .B(n3311), .Z(n3041) );
  ND2SVTX2 U1209 ( .A(n4304), .B(n4305), .Z(n4307) );
  ND2SVTX4 U1210 ( .A(n3738), .B(n3787), .Z(n3951) );
  ND3SVTX2 U1211 ( .A(n4056), .B(n3229), .C(n3230), .Z(n3228) );
  IVSVTX6 U1212 ( .A(n4056), .Z(n582) );
  AO20CSVTX4 U1213 ( .A(n3132), .B(n3179), .C(n3136), .D(n2086), .Z(n1285) );
  ND3ABSVTX4 U1214 ( .A(n3136), .B(n2082), .C(n3179), .Z(n2085) );
  IVSVTX8 U1215 ( .A(n3179), .Z(n560) );
  AO7ABSVTX6 U1216 ( .A(n633), .B(n2705), .C(n1570), .Z(n1759) );
  ND2SVTX4 U1217 ( .A(n1398), .B(n570), .Z(n3339) );
  IVSVTX8 U1218 ( .A(n376), .Z(n477) );
  AO4SVTX8 U1219 ( .A(n1072), .B(n1163), .C(n1159), .D(n1071), .Z(n1070) );
  ND2SVTX2 U1220 ( .A(n4041), .B(n4039), .Z(n4042) );
  IVSVTX12 U1221 ( .A(n1996), .Z(n2751) );
  AO7ABSVTX6 U1222 ( .A(n2579), .B(n1768), .C(n356), .Z(n2634) );
  ND2ASVTX4 U1223 ( .A(n2512), .B(n1768), .Z(n2502) );
  IVSVTX6 U1224 ( .A(n843), .Z(n2259) );
  IVSVTX2 U1225 ( .A(n4241), .Z(n4217) );
  ND2SVTX2 U1226 ( .A(n4226), .B(n1757), .Z(n4228) );
  BFSVTX10 U1227 ( .A(n4284), .Z(n339) );
  CTBUFSVTX8 U1228 ( .A(n4234), .Z(n414) );
  ENSVTX8 U1229 ( .A(n4223), .B(n4222), .Z(rslt_o[14]) );
  EOSVTX8 U1230 ( .A(n4280), .B(n4279), .Z(rslt_o[13]) );
  AO7SVTX8 U1231 ( .A(n484), .B(n366), .C(n2049), .Z(n2052) );
  AO7SVTX6 U1232 ( .A(n1465), .B(n4279), .C(n412), .Z(n4222) );
  ENSVTX8 U1233 ( .A(n1626), .B(n1624), .Z(rslt_o[17]) );
  IVSVTX4 U1234 ( .A(n3369), .Z(n568) );
  NR2ASVTX6 U1235 ( .A(n2394), .B(n1908), .Z(n4284) );
  AO6SVTX4 U1236 ( .A(n2225), .B(n4210), .C(n4209), .Z(n4211) );
  NR2ASVTX4 U1237 ( .A(n516), .B(n3215), .Z(n3321) );
  ND2ASVTX4 U1238 ( .A(n516), .B(n3215), .Z(n1491) );
  ENSVTX8 U1239 ( .A(n4193), .B(n1247), .Z(rslt_o[18]) );
  IVSVTX12 U1240 ( .A(n620), .Z(n539) );
  ND3ASVTX8 U1241 ( .A(n2421), .B(n4165), .C(n499), .Z(n4204) );
  ND4ASVTX6 U1242 ( .A(n2525), .B(n2531), .C(n2208), .D(n2228), .Z(n1147) );
  ND3SVTX2 U1243 ( .A(n3544), .B(n3545), .C(n3541), .Z(n3548) );
  ND4ASVTX4 U1244 ( .A(n1941), .B(n2561), .C(n2551), .D(n1857), .Z(n1903) );
  AN2SVTX4 U1245 ( .A(n3623), .B(n528), .Z(n2446) );
  ND2SVTX4 U1246 ( .A(n1972), .B(n1730), .Z(n3784) );
  IVSVTX6 U1247 ( .A(n2161), .Z(n559) );
  NR3SVTX6 U1248 ( .A(n4118), .B(n4119), .C(n1727), .Z(n1726) );
  CTBUFSVTX4 U1249 ( .A(n800), .Z(n366) );
  NR2ASVTX8 U1250 ( .A(n2658), .B(n1544), .Z(n1540) );
  IVSVTX12 U1251 ( .A(n2639), .Z(n632) );
  IVSVTX6 U1252 ( .A(n2582), .Z(n2503) );
  ENSVTX4 U1253 ( .A(n2885), .B(n687), .Z(n2750) );
  CTIVSVTX4 U1254 ( .A(n2237), .Z(n2015) );
  ND2SVTX8 U1255 ( .A(n2663), .B(n1974), .Z(n2125) );
  ND3SVTX8 U1256 ( .A(n2547), .B(n1108), .C(n1147), .Z(n430) );
  ND2SVTX4 U1257 ( .A(n2538), .B(n2539), .Z(n2355) );
  ND2ASVTX8 U1258 ( .A(n4001), .B(n4025), .Z(n4026) );
  AO3ABSVTX8 U1259 ( .A(n3316), .B(n1235), .C(n3313), .D(n3315), .Z(n1990) );
  ND3SVTX8 U1260 ( .A(n1990), .B(n351), .C(n1989), .Z(n1392) );
  AO7ABSVTX8 U1261 ( .A(n911), .B(n814), .C(n815), .Z(n1552) );
  IVSVTX6 U1262 ( .A(n2612), .Z(n950) );
  IVSVTX4 U1263 ( .A(n2612), .Z(n1034) );
  AO6ABSVTX4 U1264 ( .A(n3918), .B(n3920), .C(n3919), .Z(n3921) );
  BFSVTX2 U1265 ( .A(n623), .Z(n389) );
  NR3ABSVTX8 U1266 ( .A(n368), .B(n340), .C(n1775), .Z(n4268) );
  AO3SVTX6 U1267 ( .A(n1459), .B(n1463), .C(n2210), .D(n370), .Z(n340) );
  CTIVSVTX6 U1268 ( .A(n2623), .Z(n1116) );
  ND4SVTX6 U1269 ( .A(n2591), .B(n2592), .C(n2590), .D(n2576), .Z(n999) );
  ND2SVTX4 U1270 ( .A(n1576), .B(n341), .Z(n2590) );
  ND2ASVTX8 U1271 ( .A(n1921), .B(n1335), .Z(n3865) );
  IVSVTX8 U1272 ( .A(n666), .Z(n673) );
  CTIVSVTX12 U1273 ( .A(n1043), .Z(n1026) );
  ND2SVTX8 U1274 ( .A(n1119), .B(n1120), .Z(n1002) );
  IVSVTX6 U1275 ( .A(n636), .Z(n2519) );
  BFSVTX1 U1276 ( .A(num_i[5]), .Z(n343) );
  AO7SVTX8 U1277 ( .A(n2491), .B(n2552), .C(n470), .Z(n2557) );
  CTBUFSVTX8 U1278 ( .A(n1410), .Z(n861) );
  BFSVTX10 U1279 ( .A(n2678), .Z(n970) );
  ND3SVTX8 U1280 ( .A(n345), .B(n344), .C(n983), .Z(n953) );
  ND2SVTX4 U1281 ( .A(n1918), .B(n982), .Z(n344) );
  NR2SVTX4 U1282 ( .A(n987), .B(n985), .Z(n345) );
  NR2SVTX4 U1283 ( .A(n1690), .B(n1310), .Z(n1309) );
  ND3SVTX6 U1284 ( .A(n3880), .B(n1314), .C(n1312), .Z(n1310) );
  AO4SVTX6 U1285 ( .A(n1274), .B(n1273), .C(n1272), .D(n338), .Z(n2603) );
  AO7SVTX8 U1286 ( .A(n2633), .B(n1971), .C(n521), .Z(n2648) );
  NR2SVTX4 U1287 ( .A(n3866), .B(n346), .Z(n1313) );
  ND4ABSVTX8 U1288 ( .A(n347), .B(n1949), .C(n864), .D(n1948), .Z(n1084) );
  NR2SVTX4 U1289 ( .A(n3514), .B(n1343), .Z(n347) );
  ND2SVTX4 U1290 ( .A(n1576), .B(n1039), .Z(n2614) );
  AO7SVTX6 U1291 ( .A(n349), .B(n348), .C(n1791), .Z(n2060) );
  IVSVTX4 U1292 ( .A(n1330), .Z(n348) );
  IVSVTX4 U1293 ( .A(n537), .Z(n349) );
  NR2SVTX4 U1294 ( .A(n1850), .B(n569), .Z(n1503) );
  MUX21SVTX4 U1295 ( .A(n3424), .B(n3427), .S(n3426), .Z(n465) );
  BFSVTX8 U1296 ( .A(num_i[15]), .Z(n393) );
  NR2SVTX2 U1297 ( .A(n393), .B(n1755), .Z(n2468) );
  ND2SVTX4 U1298 ( .A(n1235), .B(n3317), .Z(n351) );
  AO7ASVTX8 U1299 ( .A(n3790), .B(n352), .C(n1422), .Z(n3794) );
  IVSVTX4 U1300 ( .A(n2202), .Z(n352) );
  BFSVTX12 U1301 ( .A(n501), .Z(n2017) );
  IVSVTX10 U1302 ( .A(n2308), .Z(n2126) );
  IVSVTX6 U1303 ( .A(n545), .Z(n3283) );
  EO3SVTX8 U1304 ( .A(n1268), .B(n3279), .C(n808), .Z(n2999) );
  AO4SVTX6 U1305 ( .A(n2639), .B(n970), .C(n706), .D(n820), .Z(n3279) );
  IVSVTX10 U1306 ( .A(n501), .Z(n1006) );
  AO7SVTX6 U1307 ( .A(n879), .B(n1223), .C(n1848), .Z(n1739) );
  IVSVTX10 U1308 ( .A(num_i[29]), .Z(n2486) );
  ND2SVTX6 U1309 ( .A(n690), .B(n992), .Z(n882) );
  BFSVTX8 U1310 ( .A(num_i[20]), .Z(n2534) );
  ND2SVTX8 U1311 ( .A(n1762), .B(n1323), .Z(n2670) );
  IVSVTX8 U1312 ( .A(n1124), .Z(n1115) );
  ND3SVTX8 U1313 ( .A(n1558), .B(n2378), .C(n2054), .Z(n1555) );
  IVSVTX12 U1314 ( .A(n1359), .Z(n1297) );
  AN3SVTX6 U1315 ( .A(n2424), .B(n3796), .C(n3726), .Z(n3721) );
  AO7SVTX6 U1316 ( .A(n2558), .B(n2559), .C(n2751), .Z(n949) );
  IVSVTX8 U1317 ( .A(n1967), .Z(n2849) );
  NR2ASVTX6 U1318 ( .A(n1343), .B(n3905), .Z(n2252) );
  ND2ASVTX8 U1319 ( .A(n2678), .B(n354), .Z(n1200) );
  AO4SVTX6 U1320 ( .A(n1996), .B(n2676), .C(n738), .D(n2677), .Z(n354) );
  IVSVTX8 U1321 ( .A(n1906), .Z(n1535) );
  ND3SVTX6 U1322 ( .A(n1134), .B(n355), .C(n1129), .Z(n1136) );
  ND2SVTX4 U1323 ( .A(n1133), .B(n1131), .Z(n355) );
  IVSVTX6 U1324 ( .A(n3530), .Z(n745) );
  ND3ABSVTX6 U1325 ( .A(n2671), .B(n2570), .C(n1197), .Z(n356) );
  IVSVTX4 U1326 ( .A(n796), .Z(n1852) );
  ND2ASVTX8 U1327 ( .A(n686), .B(n1058), .Z(n357) );
  NR3SVTX8 U1328 ( .A(n1785), .B(n3779), .C(n1594), .Z(n1593) );
  ND4ABSVTX8 U1329 ( .A(n3624), .B(n3866), .C(n3963), .D(n1593), .Z(n1296) );
  EO3SVTX8 U1330 ( .A(n537), .B(n2820), .C(n2819), .Z(n2823) );
  AO5ASVTX8 U1331 ( .B(n1339), .A(n1770), .C(n620), .Z(n2820) );
  ND2SVTX4 U1332 ( .A(n358), .B(n1146), .Z(n1144) );
  NR2SVTX4 U1333 ( .A(n510), .B(n3487), .Z(n358) );
  AO7ABSVTX8 U1334 ( .A(n359), .B(n500), .C(n1361), .Z(n1537) );
  IVSVTX4 U1335 ( .A(n4190), .Z(n931) );
  ND4ABSVTX8 U1336 ( .A(n1407), .B(n1262), .C(n933), .D(n934), .Z(n4190) );
  AO7SVTX6 U1337 ( .A(n3349), .B(n3350), .C(n3348), .Z(n2275) );
  ND2SVTX4 U1338 ( .A(n361), .B(n360), .Z(n1955) );
  NR2ASVTX6 U1339 ( .A(n900), .B(n2059), .Z(n360) );
  IVSVTX4 U1340 ( .A(n693), .Z(n361) );
  ND3ABSVTX4 U1341 ( .A(n1107), .B(n1061), .C(n2110), .Z(n2566) );
  NR2ASVTX6 U1342 ( .A(n2519), .B(n2585), .Z(n2542) );
  IVSVTX8 U1343 ( .A(n500), .Z(n502) );
  IVSVTX10 U1344 ( .A(n500), .Z(n503) );
  ND3SVTX8 U1345 ( .A(n1101), .B(n721), .C(n2249), .Z(n4247) );
  IVSVTX4 U1346 ( .A(n2244), .Z(n362) );
  AO6SVTX8 U1347 ( .A(n362), .B(n713), .C(n752), .Z(n3573) );
  ND2SVTX8 U1348 ( .A(n2509), .B(n2528), .Z(n1209) );
  ND2ASVTX8 U1349 ( .A(n3470), .B(n1101), .Z(n719) );
  NR2SVTX4 U1350 ( .A(n1329), .B(n1676), .Z(n3146) );
  IVSVTX4 U1351 ( .A(n454), .Z(n363) );
  ND2ASVTX8 U1352 ( .A(n363), .B(n4085), .Z(n1371) );
  AO4SVTX8 U1353 ( .A(n2598), .B(n364), .C(n786), .D(n2596), .Z(n1732) );
  ND3SVTX8 U1354 ( .A(n2593), .B(n631), .C(n2592), .Z(n364) );
  ND2SVTX4 U1355 ( .A(n1789), .B(n365), .Z(n2215) );
  ND2SVTX4 U1356 ( .A(n1790), .B(n624), .Z(n365) );
  ND3SVTX8 U1357 ( .A(n690), .B(n1108), .C(n1147), .Z(n2533) );
  IVSVTX10 U1358 ( .A(n1124), .Z(n1287) );
  EN3SVTX8 U1359 ( .A(n545), .B(n1748), .C(n808), .Z(n3070) );
  IVSVTX4 U1360 ( .A(n3070), .Z(n1370) );
  IVSVTX4 U1361 ( .A(n4247), .Z(n720) );
  IVSVTX2 U1362 ( .A(n3531), .Z(n574) );
  ND2ASVTX8 U1363 ( .A(n3531), .B(n1387), .Z(n1986) );
  ND2ASVTX8 U1364 ( .A(n3907), .B(n3492), .Z(n4249) );
  IVSVTX4 U1365 ( .A(n442), .Z(n370) );
  AO7ASVTX8 U1366 ( .A(n3453), .B(n1623), .C(n3505), .Z(n3454) );
  ND4SVTX6 U1367 ( .A(n4171), .B(n2063), .C(n848), .D(n2062), .Z(n1105) );
  IVSVTX6 U1368 ( .A(n3458), .Z(n807) );
  NR3ABSVTX8 U1369 ( .A(n3458), .B(n1551), .C(n3084), .Z(n3085) );
  IVSVTX4 U1370 ( .A(n371), .Z(n2435) );
  ND2SVTX4 U1371 ( .A(n2155), .B(n372), .Z(n371) );
  ND2SVTX4 U1372 ( .A(n2654), .B(n2587), .Z(n372) );
  IVSVTX12 U1373 ( .A(n1685), .Z(n1121) );
  IVSVTX8 U1374 ( .A(n1685), .Z(n2176) );
  BFSVTX12 U1375 ( .A(n1647), .Z(n823) );
  IVSVTX4 U1376 ( .A(n3399), .Z(n3400) );
  EO3SVTX8 U1377 ( .A(n503), .B(n617), .C(n2807), .Z(n2907) );
  ND2SVTX4 U1378 ( .A(n3282), .B(n1121), .Z(n2836) );
  IVSVTX8 U1379 ( .A(n3850), .Z(n1322) );
  IVSVTX6 U1380 ( .A(n545), .Z(n911) );
  ND2SVTX6 U1381 ( .A(n1766), .B(n3483), .Z(n2008) );
  IVSVTX8 U1382 ( .A(n2838), .Z(n2335) );
  NR3SVTX6 U1383 ( .A(n1319), .B(n930), .C(n859), .Z(n1301) );
  F_ENSVTX2 U1384 ( .A(n684), .B(n2984), .Z(n2986) );
  ND3ABSVTX8 U1385 ( .A(n1501), .B(n375), .C(n1234), .Z(n1908) );
  AO7SVTX6 U1386 ( .A(n1170), .B(n3366), .C(n3301), .Z(n376) );
  ND2SVTX4 U1387 ( .A(n377), .B(n1046), .Z(n1451) );
  ND3SVTX6 U1388 ( .A(n1454), .B(n1453), .C(n1455), .Z(n377) );
  ND3SVTX8 U1389 ( .A(n2658), .B(n1769), .C(n2232), .Z(n2541) );
  IVSVTX12 U1390 ( .A(n944), .Z(n1295) );
  IVSVTX4 U1391 ( .A(n2077), .Z(n387) );
  IVSVTX10 U1392 ( .A(n1166), .Z(n2902) );
  AO6CSVTX8 U1393 ( .A(n1981), .B(n469), .C(n2421), .Z(n4271) );
  BFSVTX8 U1394 ( .A(n1021), .Z(n648) );
  AN2SVTX8 U1395 ( .A(n2364), .B(n725), .Z(n2585) );
  ND4SVTX8 U1396 ( .A(n2220), .B(n2500), .C(n2486), .D(n2313), .Z(n666) );
  AO2SVTX6 U1397 ( .A(n2335), .B(n1052), .C(n2753), .D(n2839), .Z(n1050) );
  AO7SVTX8 U1398 ( .A(n2752), .B(n1051), .C(n1050), .Z(n2831) );
  MUX21NSVTX6 U1399 ( .A(n1308), .B(n1310), .S(n1307), .Z(n1306) );
  ND3SVTX8 U1400 ( .A(n1109), .B(n1110), .C(n379), .Z(n1533) );
  AO1SVTX8 U1401 ( .A(n698), .B(n2292), .C(n701), .D(n696), .Z(n379) );
  AO7SVTX8 U1402 ( .A(n2678), .B(n2334), .C(n380), .Z(n899) );
  ND3SVTX8 U1403 ( .A(n900), .B(n2643), .C(n2070), .Z(n380) );
  EN3SVTX8 U1404 ( .A(n1889), .B(n3068), .C(n503), .Z(n2974) );
  IVSVTX4 U1405 ( .A(n593), .Z(n3624) );
  IVSVTX4 U1406 ( .A(n381), .Z(n485) );
  ND3SVTX6 U1407 ( .A(n3583), .B(n593), .C(n3626), .Z(n381) );
  ND2ASVTX8 U1408 ( .A(n1771), .B(n382), .Z(n593) );
  IVSVTX4 U1409 ( .A(n1979), .Z(n382) );
  BFSVTX1 U1410 ( .A(n970), .Z(rslt_o[27]) );
  IVSVTX4 U1411 ( .A(n384), .Z(n761) );
  ND2SVTX4 U1412 ( .A(n1945), .B(n2714), .Z(n384) );
  AO4SVTX6 U1413 ( .A(n971), .B(n633), .C(n970), .D(n632), .Z(n1267) );
  ND4ABSVTX8 U1414 ( .A(n630), .B(n2353), .C(n385), .D(n538), .Z(n2342) );
  NR3SVTX8 U1415 ( .A(n1748), .B(n684), .C(n1647), .Z(n385) );
  IVSVTX8 U1416 ( .A(n1810), .Z(n2402) );
  ND3ABSVTX8 U1417 ( .A(n386), .B(n1898), .C(n747), .Z(n1707) );
  IVSVTX4 U1418 ( .A(n749), .Z(n386) );
  NR2SVTX8 U1419 ( .A(n1087), .B(n3442), .Z(n3526) );
  ND2SVTX6 U1420 ( .A(n970), .B(n2639), .Z(n2640) );
  ND2SVTX8 U1421 ( .A(n2442), .B(n3203), .Z(n4179) );
  BFSVTX12 U1422 ( .A(n2737), .Z(n1764) );
  ND2ASVTX8 U1423 ( .A(n1225), .B(n1743), .Z(n1224) );
  IVSVTX8 U1424 ( .A(n2308), .Z(n1768) );
  IVSVTX6 U1425 ( .A(n2353), .Z(n822) );
  BFSVTX12 U1426 ( .A(n2503), .Z(rslt_o[31]) );
  AO7ASVTX8 U1427 ( .A(n389), .B(n3923), .C(n1902), .Z(n2172) );
  IVSVTX6 U1428 ( .A(n3529), .Z(n504) );
  ND3SVTX8 U1429 ( .A(n2259), .B(n2351), .C(n2291), .Z(n3529) );
  IVSVTX8 U1430 ( .A(n3589), .Z(n1699) );
  IVSVTX12 U1431 ( .A(n1538), .Z(n1060) );
  NR2ASVTX6 U1432 ( .A(n592), .B(n3859), .Z(n3863) );
  ND2SVTX4 U1433 ( .A(n3653), .B(n3660), .Z(n3446) );
  ND3SVTX8 U1434 ( .A(n691), .B(n2264), .C(n3079), .Z(n391) );
  ND2ASVTX8 U1435 ( .A(n874), .B(n2721), .Z(n2708) );
  AO7ABSVTX8 U1436 ( .A(n2573), .B(n1756), .C(n1610), .Z(n664) );
  IVSVTX4 U1437 ( .A(n1973), .Z(n1975) );
  CTIVSVTX8 U1438 ( .A(n3564), .Z(n758) );
  BFSVTX8 U1439 ( .A(n2423), .Z(n744) );
  IVSVTX8 U1440 ( .A(n2582), .Z(n2232) );
  IVSVTX4 U1441 ( .A(n394), .Z(n3741) );
  ND2SVTX4 U1442 ( .A(n3743), .B(n3740), .Z(n394) );
  IVSVTX4 U1443 ( .A(n395), .Z(n3738) );
  NR2SVTX4 U1444 ( .A(n3096), .B(n3097), .Z(n395) );
  ND3SVTX8 U1445 ( .A(n3404), .B(n3403), .C(n1235), .Z(n3405) );
  ENSVTX6 U1446 ( .A(n2971), .B(n2150), .Z(n3606) );
  IVSVTX4 U1447 ( .A(n397), .Z(n1183) );
  AO7ABSVTX4 U1448 ( .A(n728), .B(n2905), .C(n398), .Z(n2918) );
  EO3SVTX8 U1449 ( .A(n728), .B(n2905), .C(n503), .Z(n2915) );
  ND3ABSVTX8 U1450 ( .A(n2395), .B(n521), .C(n1228), .Z(n988) );
  CTBUFSVTX8 U1451 ( .A(n1112), .Z(n1336) );
  ND2SVTX4 U1452 ( .A(n399), .B(n1121), .Z(n2837) );
  AO7SVTX8 U1453 ( .A(n411), .B(n730), .C(n2112), .Z(n2848) );
  IVSVTX12 U1454 ( .A(n1397), .Z(n2149) );
  IVSVTX12 U1455 ( .A(n1851), .Z(n2814) );
  ND3ABSVTX8 U1456 ( .A(n3141), .B(n1255), .C(n1505), .Z(n1281) );
  IVSVTX4 U1457 ( .A(n2198), .Z(n3923) );
  EO3SVTX8 U1458 ( .A(n2816), .B(n400), .C(n1801), .Z(n2198) );
  IVSVTX4 U1459 ( .A(n2815), .Z(n400) );
  IVSVTX6 U1460 ( .A(n646), .Z(n795) );
  IVSVTX12 U1461 ( .A(n795), .Z(n512) );
  IVSVTX4 U1462 ( .A(n2853), .Z(n2857) );
  AO7SVTX8 U1463 ( .A(n2857), .B(n1912), .C(n2856), .Z(n2237) );
  AO21SVTX8 U1464 ( .A(n404), .B(n488), .C(n3467), .D(n2251), .Z(n2250) );
  IVSVTX4 U1465 ( .A(n406), .Z(n405) );
  NR2SVTX4 U1466 ( .A(n3465), .B(n577), .Z(n406) );
  AO7ABSVTX6 U1467 ( .A(n1892), .B(n814), .C(n2977), .Z(n2980) );
  AO17SVTX8 U1468 ( .A(n1205), .B(n3857), .C(n3418), .D(n1203), .Z(n3235) );
  IVSVTX4 U1469 ( .A(n407), .Z(n2145) );
  ND2SVTX4 U1470 ( .A(num_i[1]), .B(n2507), .Z(n407) );
  EO3SVTX8 U1471 ( .A(n1889), .B(n3280), .C(n942), .Z(n2919) );
  IVSVTX8 U1472 ( .A(n2514), .Z(n1239) );
  IVSVTX12 U1473 ( .A(n1538), .Z(n1323) );
  BFSVTX4 U1474 ( .A(n1085), .Z(n408) );
  ND2SVTX8 U1475 ( .A(n3651), .B(n3652), .Z(n1832) );
  ND2ASVTX8 U1476 ( .A(n410), .B(n1539), .Z(n827) );
  IVSVTX8 U1477 ( .A(n3311), .Z(n609) );
  IVSVTX4 U1478 ( .A(n1199), .Z(n411) );
  BFSVTX1 U1479 ( .A(n4278), .Z(n412) );
  IVSVTX12 U1480 ( .A(n3654), .Z(n2424) );
  ND2SVTX4 U1481 ( .A(n707), .B(n649), .Z(n952) );
  AO7SVTX8 U1482 ( .A(n3501), .B(n1128), .C(n3502), .Z(n3456) );
  ND2SVTX4 U1483 ( .A(n2243), .B(n1094), .Z(n2415) );
  ND2SVTX4 U1484 ( .A(n417), .B(n416), .Z(n634) );
  IVSVTX4 U1485 ( .A(n2581), .Z(n417) );
  AO7SVTX8 U1486 ( .A(n1365), .B(n477), .C(n419), .Z(n1269) );
  AO6SVTX8 U1487 ( .A(n582), .B(n581), .C(n580), .Z(n419) );
  NR2SVTX4 U1488 ( .A(n1381), .B(n420), .Z(n1380) );
  ND3SVTX6 U1489 ( .A(n1385), .B(n2241), .C(n421), .Z(n420) );
  AO7SVTX6 U1490 ( .A(n1383), .B(n1384), .C(n4066), .Z(n421) );
  ND3SVTX6 U1491 ( .A(n1824), .B(n423), .C(n422), .Z(n1821) );
  IVSVTX4 U1492 ( .A(n3710), .Z(n423) );
  ENSVTX8 U1493 ( .A(n424), .B(n2417), .Z(n4133) );
  ENSVTX8 U1494 ( .A(n2794), .B(n591), .Z(n424) );
  NR2SVTX4 U1495 ( .A(n426), .B(n425), .Z(n2094) );
  IVSVTX4 U1496 ( .A(n2099), .Z(n425) );
  AO6SVTX4 U1497 ( .A(n3265), .B(n3266), .C(n2381), .Z(n426) );
  IVSVTX10 U1498 ( .A(n900), .Z(n1043) );
  IVSVTX6 U1499 ( .A(n2849), .Z(n2137) );
  IVSVTX12 U1500 ( .A(n1090), .Z(n1647) );
  IVSVTX6 U1501 ( .A(n2751), .Z(n2306) );
  BFSVTX1 U1502 ( .A(n4258), .Z(n429) );
  IVSVTX10 U1503 ( .A(n1023), .Z(n1022) );
  IVSVTX4 U1504 ( .A(n430), .Z(n471) );
  ND3SVTX8 U1505 ( .A(n2067), .B(n731), .C(n2074), .Z(n2072) );
  AO7SVTX8 U1506 ( .A(n2072), .B(n852), .C(n2071), .Z(n2106) );
  AO6SVTX8 U1507 ( .A(n2100), .B(n2807), .C(n2743), .Z(n2714) );
  AO4SVTX8 U1508 ( .A(n2834), .B(n2835), .C(n3067), .D(n2833), .Z(n1024) );
  ND2ASVTX8 U1509 ( .A(n4073), .B(n781), .Z(n2382) );
  IVSVTX8 U1510 ( .A(num_i[25]), .Z(n637) );
  AO6SVTX4 U1511 ( .A(n1036), .B(n2503), .C(n2553), .Z(n2556) );
  NR2ASVTX6 U1512 ( .A(n2584), .B(n431), .Z(n2333) );
  ND2ASVTX8 U1513 ( .A(n3079), .B(n3075), .Z(n3505) );
  BFSVTX6 U1514 ( .A(n4058), .Z(n433) );
  NR2SVTX4 U1515 ( .A(n3432), .B(n1963), .Z(n1958) );
  ND2SVTX4 U1516 ( .A(n3288), .B(n434), .Z(n3432) );
  IVSVTX4 U1517 ( .A(n614), .Z(n434) );
  ND2SVTX4 U1518 ( .A(n2887), .B(n687), .Z(n3477) );
  IVSVTX8 U1519 ( .A(n1541), .Z(n2680) );
  AO2ABSVTX4 U1520 ( .C(n3076), .D(n3075), .A(n3074), .B(n3079), .Z(n3077) );
  ND3SVTX8 U1521 ( .A(n3448), .B(n3447), .C(n2436), .Z(n1101) );
  NR3SVTX8 U1522 ( .A(n438), .B(n2516), .C(n2515), .Z(n2476) );
  NR3SVTX8 U1523 ( .A(num_i[10]), .B(num_i[11]), .C(n2472), .Z(n438) );
  BFSVTX12 U1524 ( .A(n1361), .Z(n1223) );
  IVSVTX4 U1525 ( .A(n2000), .Z(n1999) );
  ND3SVTX8 U1526 ( .A(n1999), .B(n1998), .C(n2001), .Z(n3234) );
  IVSVTX6 U1527 ( .A(n2552), .Z(n654) );
  IVSVTX12 U1528 ( .A(n2570), .Z(n2308) );
  IVSVTX2 U1529 ( .A(n880), .Z(n1133) );
  EO3SVTX8 U1530 ( .A(n798), .B(n686), .C(n3078), .Z(n3081) );
  IVSVTX8 U1531 ( .A(n1643), .Z(n661) );
  IVSVTX4 U1532 ( .A(n440), .Z(n1868) );
  ND2SVTX4 U1533 ( .A(n2724), .B(n2725), .Z(n440) );
  IVSVTX6 U1534 ( .A(n1117), .Z(n1112) );
  ND2ASVTX8 U1535 ( .A(n2973), .B(n2300), .Z(n3625) );
  ND3SVTX8 U1536 ( .A(n746), .B(n556), .C(n1202), .Z(n4205) );
  AO21SVTX8 U1537 ( .A(n3156), .B(n3153), .C(n960), .D(n561), .Z(n3149) );
  ND3ABSVTX8 U1538 ( .A(n4073), .B(n3119), .C(n3120), .Z(n442) );
  IVSVTX8 U1539 ( .A(n1021), .Z(n878) );
  AO4ABSVTX6 U1540 ( .C(n670), .D(n878), .A(n668), .B(n761), .Z(n696) );
  IVSVTX6 U1541 ( .A(n1118), .Z(n2243) );
  IVSVTX10 U1542 ( .A(n2243), .Z(n2612) );
  AO7SVTX8 U1543 ( .A(n2483), .B(n1341), .C(n1744), .Z(n2484) );
  IVSVTX12 U1544 ( .A(n1346), .Z(n616) );
  AO7CSVTX6 U1545 ( .A(n1361), .B(n541), .C(n616), .Z(n1362) );
  ND2SVTX4 U1546 ( .A(n4206), .B(n4204), .Z(n4208) );
  IVSVTX8 U1547 ( .A(n3396), .Z(n3055) );
  NR3ABSVTX8 U1548 ( .A(n2255), .B(n2784), .C(n443), .Z(n2709) );
  IVSVTX4 U1549 ( .A(n542), .Z(n443) );
  ND2ASVTX8 U1550 ( .A(n1600), .B(n1745), .Z(n2804) );
  IVSVTX10 U1551 ( .A(n3260), .Z(n558) );
  ND4SVTX6 U1552 ( .A(n1388), .B(n2498), .C(n2377), .D(n2492), .Z(n1682) );
  AO6SVTX4 U1553 ( .A(n3882), .B(n447), .C(n3686), .Z(n446) );
  NR2SVTX4 U1554 ( .A(n2399), .B(n1690), .Z(n447) );
  ND2ASVTX8 U1555 ( .A(n1823), .B(n812), .Z(n3772) );
  AO17SVTX4 U1556 ( .A(n3450), .B(n2884), .C(n2886), .D(n3508), .Z(n832) );
  ND2ASVTX8 U1557 ( .A(n448), .B(n2316), .Z(n3508) );
  IVSVTX4 U1558 ( .A(n517), .Z(n448) );
  IVSVTX4 U1559 ( .A(n2626), .Z(n676) );
  ND4ABSVTX8 U1560 ( .A(n3869), .B(n3868), .C(n2118), .D(n1322), .Z(n3906) );
  NR3SVTX8 U1561 ( .A(n3864), .B(n3863), .C(n3862), .Z(n3869) );
  IVSVTX8 U1562 ( .A(num_i[26]), .Z(n640) );
  IVSVTX8 U1563 ( .A(n2801), .Z(n771) );
  BFSVTX1 U1564 ( .A(n647), .Z(n450) );
  BFSVTX1 U1565 ( .A(num_i[4]), .Z(n451) );
  AO7ABSVTX8 U1566 ( .A(n2036), .B(n2183), .C(n2616), .Z(n1152) );
  ND3SVTX8 U1567 ( .A(n2715), .B(n695), .C(n3241), .Z(n694) );
  ND3SVTX8 U1568 ( .A(n2142), .B(n2288), .C(n2714), .Z(n3241) );
  IVSVTX8 U1569 ( .A(n664), .Z(n2184) );
  IVSVTX4 U1570 ( .A(n723), .Z(n722) );
  NR3ABSVTX8 U1571 ( .A(n1182), .B(n452), .C(n1180), .Z(n1188) );
  ND3ASVTX6 U1572 ( .A(n3954), .B(n1879), .C(n3953), .Z(n452) );
  ND2ASVTX8 U1573 ( .A(n3856), .B(n3855), .Z(n3859) );
  EO3SVTX8 U1574 ( .A(n2398), .B(n539), .C(n2868), .Z(n2773) );
  AO7SVTX8 U1575 ( .A(n2775), .B(n3382), .C(n3352), .Z(n2350) );
  NR2SVTX2 U1576 ( .A(n428), .B(n2883), .Z(n688) );
  ND3SVTX4 U1577 ( .A(n949), .B(n680), .C(n2560), .Z(n947) );
  IVSVTX4 U1578 ( .A(n2618), .Z(n1576) );
  IVSVTX0H U1579 ( .A(n2982), .Z(n2983) );
  F_ND2ASVTX2 U1580 ( .A(n2081), .B(n2636), .Z(n2575) );
  NR2SVTX2 U1581 ( .A(n546), .B(n2858), .Z(n2051) );
  CTBUFSVTX12 U1582 ( .A(n519), .Z(n1518) );
  IVSVTX2 U1583 ( .A(n3054), .Z(n1985) );
  F_ND2ASVTX2 U1584 ( .A(n4120), .B(n4121), .Z(n1727) );
  F_ND3SVTX2 U1585 ( .A(n2067), .B(n3969), .C(n3970), .Z(n3971) );
  NR2SVTX0H U1586 ( .A(n3384), .B(n3362), .Z(n3361) );
  F_AN2SVTX2 U1587 ( .A(n3111), .B(n606), .Z(n2412) );
  ND2SVTX2 U1588 ( .A(n485), .B(n3865), .Z(n1307) );
  ND2SVTX4 U1589 ( .A(n3744), .B(n1729), .Z(n3757) );
  IVSVTX2 U1590 ( .A(n638), .Z(n2513) );
  F_ND2ASVTX2 U1591 ( .A(n538), .B(n2352), .Z(n1951) );
  BFSVTX2 U1592 ( .A(n1796), .Z(n1636) );
  IVSVTX4 U1593 ( .A(n3613), .Z(n1343) );
  BFSVTX0H U1594 ( .A(n4050), .Z(n4051) );
  IVSVTX0H U1595 ( .A(n4176), .Z(n597) );
  AO6SVTX1 U1596 ( .A(n4181), .B(n2303), .C(n1660), .Z(n2302) );
  ND3SVTX4 U1597 ( .A(n2467), .B(n2298), .C(n1806), .Z(n973) );
  IVSVTX0H U1598 ( .A(n2421), .Z(n4149) );
  IVSVTX0H U1599 ( .A(n1866), .Z(n2766) );
  F_AN2SVTX2 U1600 ( .A(n1596), .B(n4074), .Z(n454) );
  F_EOSVTX2 U1601 ( .A(n2985), .B(n2765), .Z(n455) );
  F_EOSVTX2 U1602 ( .A(n3441), .B(n2755), .Z(n457) );
  AO7NSVTX2 U1603 ( .A(n4159), .B(n739), .C(n594), .Z(n458) );
  OR2SVTX4 U1604 ( .A(n1223), .B(n623), .Z(n459) );
  F_AN2SVTX2 U1605 ( .A(n3829), .B(n3834), .Z(n461) );
  AN2SVTX4 U1606 ( .A(n3851), .B(n2455), .Z(n462) );
  AN2SVTX4 U1607 ( .A(n1937), .B(n643), .Z(n463) );
  AO7NSVTX4 U1608 ( .A(n3945), .B(n3944), .C(n1340), .Z(n464) );
  BFSVTX6 U1609 ( .A(num_i[17]), .Z(n892) );
  F_AN2SVTX2 U1610 ( .A(n4174), .B(n2350), .Z(n467) );
  F_MUX21SVTX2 U1611 ( .A(n3704), .B(n1040), .S(n3712), .Z(n468) );
  AO7NSVTX6 U1612 ( .A(n4085), .B(n4084), .C(n4083), .Z(n469) );
  AN2SVTX4 U1613 ( .A(n920), .B(n2582), .Z(n470) );
  IVSVTX8 U1614 ( .A(n2678), .Z(n820) );
  IVSVTX10 U1615 ( .A(n1083), .Z(n633) );
  IVSVTX12 U1616 ( .A(n1359), .Z(n1360) );
  CTOR3SVTX4 U1617 ( .A(n2628), .B(n1701), .C(n738), .Z(n472) );
  IVSVTX10 U1618 ( .A(n1323), .Z(n1996) );
  IVSVTX12 U1619 ( .A(n2905), .Z(n623) );
  AN2SVTX4 U1620 ( .A(n1939), .B(n1481), .Z(n473) );
  CTBUFSVTX8 U1621 ( .A(n1939), .Z(n964) );
  ND2SVTX2 U1622 ( .A(n1717), .B(n619), .Z(n824) );
  IVSVTX8 U1623 ( .A(n1536), .Z(n2865) );
  IVSVTX10 U1624 ( .A(n1642), .Z(n2344) );
  NR2ASVTX2 U1625 ( .A(n2760), .B(n3283), .Z(n729) );
  AO7SVTX8 U1626 ( .A(n3441), .B(n3440), .C(n3439), .Z(n1662) );
  IVSVTX8 U1627 ( .A(n1662), .Z(n2420) );
  IVSVTX10 U1628 ( .A(n1546), .Z(n1547) );
  ND2ASVTX8 U1629 ( .A(n3111), .B(n4133), .Z(n1494) );
  ND2SVTX2 U1630 ( .A(n3036), .B(n3035), .Z(n4150) );
  F_EOSVTX2 U1631 ( .A(n2759), .B(n3453), .Z(n474) );
  F_EOSVTX2 U1632 ( .A(n3436), .B(n2034), .Z(n475) );
  F_EOSVTX2 U1633 ( .A(n3521), .B(n3520), .Z(n476) );
  F_AN2SVTX2 U1634 ( .A(n2348), .B(n1334), .Z(n478) );
  F_AN2SVTX2 U1635 ( .A(n3722), .B(n3725), .Z(n479) );
  IVSVTX2 U1636 ( .A(n1991), .Z(n2158) );
  AN2SVTX4 U1637 ( .A(n1173), .B(n1329), .Z(n480) );
  ND2ASVTX8 U1638 ( .A(n2462), .B(n2771), .Z(n2772) );
  AO5ASVTX6 U1639 ( .B(n2223), .A(n1764), .C(n3270), .Z(n1907) );
  AN2SVTX4 U1640 ( .A(n3933), .B(n3393), .Z(n482) );
  AN2SVTX4 U1641 ( .A(n3377), .B(n509), .Z(n483) );
  CTBUFSVTX8 U1642 ( .A(n2374), .Z(n974) );
  AN3SVTX8 U1643 ( .A(n1303), .B(n1302), .C(n1301), .Z(n486) );
  AO7SVTX8 U1644 ( .A(n3926), .B(n3925), .C(n3924), .Z(n3995) );
  IVSVTX6 U1645 ( .A(n3995), .Z(n3996) );
  ND2ASVTX8 U1646 ( .A(n2979), .B(n2189), .Z(n2190) );
  F_EOSVTX2 U1647 ( .A(n3488), .B(n1824), .Z(n487) );
  AN2SVTX4 U1648 ( .A(n3473), .B(n3469), .Z(n488) );
  IVSVTX4 U1649 ( .A(n3873), .Z(n928) );
  ND2SVTX4 U1650 ( .A(n2904), .B(n2903), .Z(n3852) );
  IVSVTX4 U1651 ( .A(n1739), .Z(n3060) );
  AN3SVTX4 U1652 ( .A(n1328), .B(n793), .C(n570), .Z(n489) );
  IVSVTX4 U1653 ( .A(n679), .Z(n3986) );
  AO4NSVTX4 U1654 ( .A(n3957), .B(n3959), .C(n3958), .D(n1921), .Z(n491) );
  IVSVTX4 U1655 ( .A(n1313), .Z(n1312) );
  AN2SVTX4 U1656 ( .A(n1669), .B(n962), .Z(n492) );
  AN3SVTX6 U1657 ( .A(n3790), .B(n3929), .C(n1864), .Z(n494) );
  IVSVTX10 U1658 ( .A(n1777), .Z(n765) );
  AN2SVTX4 U1659 ( .A(n2971), .B(n1777), .Z(n495) );
  AO6NSVTX4 U1660 ( .A(n2210), .B(n3120), .C(n3116), .Z(n496) );
  ND2SVTX2 U1661 ( .A(n3119), .B(n4171), .Z(n3116) );
  NR2ASVTX1 U1662 ( .A(n3383), .B(n3528), .Z(n763) );
  IVSVTX12 U1663 ( .A(n4073), .Z(n514) );
  AO7NSVTX4 U1664 ( .A(n4069), .B(n1705), .C(n514), .Z(n497) );
  ND2SVTX4 U1665 ( .A(n514), .B(n3355), .Z(n1097) );
  ND2SVTX2 U1666 ( .A(n527), .B(n3147), .Z(n2421) );
  ND3ABSVTX2 U1667 ( .A(n3429), .B(n588), .C(n3490), .Z(n1619) );
  AO4NSVTX8 U1668 ( .A(n1446), .B(n1780), .C(n498), .D(n1781), .Z(n499) );
  AO7SVTX8 U1669 ( .A(n3993), .B(n3994), .C(n1670), .Z(n1014) );
  ENSVTX6 U1670 ( .A(n2151), .B(n1940), .Z(n2990) );
  AO6ASVTX8 U1671 ( .A(n3435), .B(n3518), .C(n3434), .Z(n3534) );
  AO1CDSVTX4 U1672 ( .A(n1235), .B(n568), .C(n3368), .D(n1422), .Z(n1241) );
  IVSVTX8 U1673 ( .A(n1977), .Z(n3897) );
  AO5ASVTX6 U1674 ( .B(n2817), .A(n610), .C(n1342), .Z(n2825) );
  F_ND2ASVTX2 U1675 ( .A(n4119), .B(n3322), .Z(n3330) );
  AO7SVTX6 U1676 ( .A(n1661), .B(n727), .C(n3457), .Z(n3072) );
  IVSVTX4 U1677 ( .A(n819), .Z(n3003) );
  IVSVTX2 U1678 ( .A(n2516), .Z(n2365) );
  NR2SVTX2 U1679 ( .A(n3416), .B(n3415), .Z(n1905) );
  AO6ABSVTX8 U1680 ( .A(n1153), .B(n1421), .C(n2608), .Z(n1155) );
  EO3SVTX6 U1681 ( .A(n1419), .B(n4018), .C(n617), .Z(n2819) );
  IVSVTX4 U1682 ( .A(n4018), .Z(n1339) );
  IVSVTX6 U1683 ( .A(n4018), .Z(n3059) );
  EO3SVTX8 U1684 ( .A(n944), .B(n1518), .C(n2807), .Z(n2185) );
  ND2SVTX4 U1685 ( .A(n2724), .B(n2725), .Z(n2100) );
  ND3SVTX4 U1686 ( .A(n2724), .B(n2725), .C(n598), .Z(n2343) );
  BFSVTX12 U1687 ( .A(n1166), .Z(n2576) );
  AO6SVTX4 U1688 ( .A(n2240), .B(n2971), .C(n519), .Z(n994) );
  IVSVTX8 U1689 ( .A(n1199), .Z(n1644) );
  IVSVTX8 U1690 ( .A(n1199), .Z(n547) );
  ND2SVTX2 U1691 ( .A(n1805), .B(n646), .Z(n645) );
  IVSVTX4 U1692 ( .A(n4204), .Z(n4166) );
  ND3SVTX8 U1693 ( .A(n2698), .B(n2245), .C(n1219), .Z(n2506) );
  IVSVTX12 U1694 ( .A(n1090), .Z(n1685) );
  AO7SVTX6 U1695 ( .A(n623), .B(n2968), .C(n2967), .Z(n3724) );
  AO7SVTX4 U1696 ( .A(n2144), .B(n861), .C(n2209), .Z(n2208) );
  ND3ABSVTX4 U1697 ( .A(n3116), .B(n3260), .C(n4167), .Z(n1469) );
  AO2SVTX4 U1698 ( .A(n1460), .B(n4091), .C(n558), .D(n4167), .Z(n1459) );
  NR2SVTX2 U1699 ( .A(n2398), .B(n1361), .Z(n1225) );
  IVSVTX8 U1700 ( .A(n2321), .Z(n835) );
  AO17CSVTX4 U1701 ( .A(n767), .B(n3018), .C(n2943), .D(n764), .Z(n1076) );
  ND2SVTX2 U1702 ( .A(n1915), .B(n3454), .Z(n3455) );
  ENSVTX6 U1703 ( .A(n777), .B(n1295), .Z(n779) );
  NR3SVTX8 U1704 ( .A(n2814), .B(n2733), .C(n2732), .Z(n2740) );
  ND2SVTX4 U1705 ( .A(n3789), .B(n3172), .Z(n4032) );
  BFSVTX8 U1706 ( .A(n3789), .Z(n1838) );
  AO7CSVTX4 U1707 ( .A(n1698), .B(n4023), .C(n2014), .Z(n4024) );
  AO2SVTX8 U1708 ( .A(n2359), .B(n2428), .C(n2286), .D(n3803), .Z(n3804) );
  IVSVTX6 U1709 ( .A(n4018), .Z(n943) );
  ND2SVTX4 U1710 ( .A(n2320), .B(n1092), .Z(n646) );
  IVSVTX12 U1711 ( .A(n3059), .Z(n500) );
  ND3ABSVTX4 U1712 ( .A(n555), .B(n2570), .C(n1197), .Z(n1672) );
  FAS1SVTX4 U1713 ( .A(n944), .B(n540), .CI(n620), .CO(n3038), .Z(n3056) );
  IVSVTX8 U1714 ( .A(n2239), .Z(n2286) );
  ND2SVTX4 U1715 ( .A(n1983), .B(n1945), .Z(n3240) );
  ND3ABSVTX6 U1716 ( .A(n2387), .B(n2727), .C(n1945), .Z(n2119) );
  ND4SVTX8 U1717 ( .A(n1210), .B(n834), .C(n1957), .D(n2656), .Z(n1954) );
  ND4SVTX8 U1718 ( .A(n2550), .B(n1083), .C(n2549), .D(n946), .Z(n945) );
  IVSVTX4 U1719 ( .A(n952), .Z(n946) );
  IVSVTX8 U1720 ( .A(n2657), .Z(n900) );
  F_EOSVTX2 U1721 ( .A(n4265), .B(n4264), .Z(rslt_o[2]) );
  AO17SVTX4 U1722 ( .A(n557), .B(n2099), .C(n2095), .D(n2093), .Z(n938) );
  AO7SVTX4 U1723 ( .A(n3407), .B(n3406), .C(n3405), .Z(n3408) );
  ND2SVTX4 U1724 ( .A(n4115), .B(n4109), .Z(n3144) );
  B_ND2SVTX2 U1725 ( .A(n1531), .B(n3225), .Z(n3226) );
  B_ND2SVTX2 U1726 ( .A(n679), .B(n736), .Z(n735) );
  ND2SVTX2 U1727 ( .A(n3988), .B(n679), .Z(n3991) );
  B_ND2SVTX2 U1728 ( .A(n4163), .B(n4162), .Z(n4164) );
  ND2SVTX2 U1729 ( .A(n3157), .B(n1430), .Z(n1429) );
  NR2SVTX2 U1730 ( .A(n1176), .B(n3987), .Z(n3988) );
  CTIVSVTX2 U1731 ( .A(n3987), .Z(n736) );
  ND2SVTX2 U1732 ( .A(n441), .B(n626), .Z(n2241) );
  B_ND2SVTX2 U1733 ( .A(n461), .B(n926), .Z(n925) );
  NR3SVTX2 U1734 ( .A(n3710), .B(n1449), .C(n576), .Z(n1448) );
  CTIVSVTX2 U1735 ( .A(n4059), .Z(n4060) );
  IVSVTX8 U1736 ( .A(n1432), .Z(n3660) );
  IVSVTX6 U1737 ( .A(n844), .Z(n583) );
  IVSVTX2 U1738 ( .A(n3765), .Z(n3767) );
  IVSVTX2 U1739 ( .A(n3998), .Z(n2809) );
  CTIVSVTX2 U1740 ( .A(n3895), .Z(n3896) );
  IVSVTX2 U1741 ( .A(n885), .Z(n2373) );
  NR2SVTX6 U1742 ( .A(n2862), .B(n2861), .Z(n1432) );
  ND2SVTX4 U1743 ( .A(n1751), .B(n2216), .Z(n4056) );
  B_ND2SVTX2 U1744 ( .A(n1790), .B(n2826), .Z(n4135) );
  ND2SVTX2 U1745 ( .A(n1482), .B(n1572), .Z(n2795) );
  CTIVSVTX2 U1746 ( .A(n505), .Z(n1508) );
  ND2SVTX2 U1747 ( .A(n2944), .B(n2865), .Z(n1572) );
  CTIVSVTX2 U1748 ( .A(n3428), .Z(n1786) );
  B_ND2SVTX2 U1749 ( .A(n506), .B(n540), .Z(n2930) );
  ND2ASVTX6 U1750 ( .A(n2893), .B(n2261), .Z(n3661) );
  CTIVSVTX2 U1751 ( .A(n516), .Z(n2940) );
  IVSVTX10 U1752 ( .A(n1547), .Z(n506) );
  ND2SVTX4 U1753 ( .A(n2893), .B(n2892), .Z(n2154) );
  IVSVTX2 U1754 ( .A(n4007), .Z(n1993) );
  NR2SVTX2 U1755 ( .A(n507), .B(n610), .Z(n1600) );
  IVSVTX2 U1756 ( .A(n2916), .Z(n1684) );
  CTIVSVTX4 U1757 ( .A(n841), .Z(n1553) );
  IVSVTX2 U1758 ( .A(n2776), .Z(n2341) );
  CTIVSVTX2 U1759 ( .A(n3495), .Z(n3515) );
  B_ND2SVTX2 U1760 ( .A(n3079), .B(n3073), .Z(n3076) );
  IVSVTX10 U1761 ( .A(n2720), .Z(n3024) );
  IVSVTX10 U1762 ( .A(n675), .Z(n3079) );
  ND2SVTX2 U1763 ( .A(n548), .B(n2983), .Z(n2984) );
  NR2SVTX2 U1764 ( .A(n2689), .B(n2685), .Z(n2683) );
  CTIVSVTX2 U1765 ( .A(n2686), .Z(n2687) );
  NR2ASVTX4 U1766 ( .A(n552), .B(n2697), .Z(n2332) );
  IVSVTX2 U1767 ( .A(n2395), .Z(n965) );
  IVSVTX2 U1768 ( .A(n1543), .Z(n1542) );
  IVSVTX10 U1769 ( .A(n2621), .Z(n2364) );
  B_ND2SVTX2 U1770 ( .A(n4294), .B(n4293), .Z(n4303) );
  ND3SVTX4 U1771 ( .A(n938), .B(n936), .C(n937), .Z(n935) );
  ENSVTX4 U1772 ( .A(n2432), .B(n4267), .Z(rslt_o[1]) );
  ND3ABSVTX4 U1773 ( .A(n2233), .B(n465), .C(n2187), .Z(n2186) );
  IVSVTX2 U1774 ( .A(n2139), .Z(n3152) );
  ND3ABSVTX4 U1775 ( .A(n1635), .B(n787), .C(n3376), .Z(n3331) );
  IVSVTX2 U1776 ( .A(n2400), .Z(n1463) );
  IVSVTX2 U1777 ( .A(n514), .Z(n1406) );
  B_ND2SVTX2 U1778 ( .A(n733), .B(n1983), .Z(n2166) );
  NR2SVTX2 U1779 ( .A(n754), .B(n3838), .Z(n3849) );
  IVSVTX4 U1780 ( .A(n4153), .Z(n525) );
  ND2SVTX2 U1781 ( .A(n3210), .B(n3208), .Z(n3207) );
  IVSVTX2 U1782 ( .A(n2097), .Z(n2096) );
  B_ND2SVTX2 U1783 ( .A(n3068), .B(n441), .Z(n2293) );
  B_ND2SVTX2 U1784 ( .A(n4100), .B(n4099), .Z(n4104) );
  CTIVSVTX2 U1785 ( .A(n3937), .Z(n3944) );
  ND2SVTX2 U1786 ( .A(n3835), .B(n3830), .Z(n927) );
  CTIVSVTX2 U1787 ( .A(n3940), .Z(n3941) );
  AN2SVTX6 U1788 ( .A(n4121), .B(n3201), .Z(n2456) );
  IVSVTX2 U1789 ( .A(n2929), .Z(n4099) );
  ND2ASVTX4 U1790 ( .A(n742), .B(n3301), .Z(n3307) );
  B_ND2SVTX2 U1791 ( .A(n3763), .B(n1884), .Z(n1883) );
  ND2SVTX2 U1792 ( .A(n589), .B(n578), .Z(n2932) );
  ND2ASVTX4 U1793 ( .A(n1409), .B(n575), .Z(n3946) );
  CTIVSVTX2 U1794 ( .A(n3709), .Z(n1449) );
  B_ND2SVTX2 U1795 ( .A(n2927), .B(n2926), .Z(n3166) );
  IVSVTX2 U1796 ( .A(n3875), .Z(n876) );
  CTIVSVTX2 U1797 ( .A(n590), .Z(n1966) );
  B_ND2SVTX2 U1798 ( .A(n3394), .B(n4030), .Z(n3395) );
  F_AN2SVTX2 U1799 ( .A(n4150), .B(n4152), .Z(n3106) );
  ND2SVTX6 U1800 ( .A(n773), .B(n774), .Z(n1719) );
  ND3SVTX4 U1801 ( .A(n3047), .B(n3390), .C(n3055), .Z(n1396) );
  NR2SVTX4 U1802 ( .A(n2979), .B(n2980), .Z(n1785) );
  IVSVTX4 U1803 ( .A(n595), .Z(n1040) );
  NR2SVTX2 U1804 ( .A(n1825), .B(n3671), .Z(n3679) );
  CTIVSVTX2 U1805 ( .A(n3487), .Z(n1816) );
  IVSVTX0H U1806 ( .A(n4120), .Z(n4116) );
  AN2SVTX6 U1807 ( .A(n3638), .B(n2347), .Z(n3889) );
  IVSVTX6 U1808 ( .A(n2154), .Z(n510) );
  ND2SVTX4 U1809 ( .A(n3024), .B(n2717), .Z(n2742) );
  B_ND2SVTX2 U1810 ( .A(n2754), .B(n3439), .Z(n2755) );
  IVSVTX6 U1811 ( .A(n3662), .Z(n505) );
  IVSVTX2 U1812 ( .A(n3010), .Z(n604) );
  IVSVTX4 U1813 ( .A(n2814), .Z(n2199) );
  IVSVTX2 U1814 ( .A(n824), .Z(n1825) );
  IVSVTX4 U1815 ( .A(n1481), .Z(n612) );
  CTBUFSVTX12 U1816 ( .A(n2398), .Z(n2807) );
  IVSVTX6 U1817 ( .A(n546), .Z(n962) );
  IVSVTX8 U1818 ( .A(n1267), .Z(n546) );
  IVSVTX12 U1819 ( .A(n3079), .Z(n508) );
  CTIVSVTX2 U1820 ( .A(n2673), .Z(n1047) );
  IVSVTX6 U1821 ( .A(n512), .Z(n521) );
  CTIVSVTX2 U1822 ( .A(n2312), .Z(n2633) );
  CTIVSVTX4 U1823 ( .A(n2365), .Z(n2366) );
  NR2SVTX2 U1824 ( .A(n555), .B(n1388), .Z(n1568) );
  ND2SVTX6 U1825 ( .A(n4290), .B(n1391), .Z(n4273) );
  NR3ABSVTX6 U1826 ( .A(n1431), .B(n4149), .C(n3200), .Z(n4196) );
  CTIVSVTX4 U1827 ( .A(n3020), .Z(n1562) );
  ND2SVTX2 U1828 ( .A(n458), .B(n2221), .Z(n1442) );
  NR4ABCSVTX4 U1829 ( .A(n3154), .B(n3156), .C(n3155), .D(n1645), .Z(n3159) );
  IVSVTX2 U1830 ( .A(n414), .Z(n4244) );
  CTIVSVTX2 U1831 ( .A(n4235), .Z(n4236) );
  CTIVSVTX2 U1832 ( .A(n2182), .Z(n2181) );
  AO8ASVTX2 U1833 ( .A(n597), .B(n4110), .C(n961), .D(n2166), .Z(n2165) );
  IVSVTX2 U1834 ( .A(n1158), .Z(n1156) );
  ND2SVTX6 U1835 ( .A(n566), .B(n954), .Z(n4235) );
  NR2SVTX2 U1836 ( .A(n4162), .B(n4155), .Z(n2221) );
  AO17SVTX2 U1837 ( .A(n3210), .B(n3209), .C(n3208), .D(n3207), .Z(n2121) );
  CTIVSVTX2 U1838 ( .A(n4063), .Z(n2091) );
  ND3ABSVTX4 U1839 ( .A(n532), .B(n3168), .C(n2362), .Z(n1505) );
  AO1CDSVTX4 U1840 ( .A(n560), .B(n4159), .C(n1931), .D(n3057), .Z(n1573) );
  ND3SVTX6 U1841 ( .A(n1103), .B(n1105), .C(n1104), .Z(n3561) );
  IVSVTX2 U1842 ( .A(n1028), .Z(n1027) );
  ND2ASVTX4 U1843 ( .A(n1777), .B(n504), .Z(n3688) );
  CTIVSVTX2 U1844 ( .A(n3355), .Z(n3354) );
  AN2SVTX6 U1845 ( .A(n589), .B(n4141), .Z(n4144) );
  ND3SVTX4 U1846 ( .A(n3996), .B(n3946), .C(n1530), .Z(n1028) );
  ND2ASVTX6 U1847 ( .A(n1293), .B(n3294), .Z(n3297) );
  CTIVSVTX4 U1848 ( .A(n2346), .Z(n3214) );
  CTIVSVTX2 U1849 ( .A(n4104), .Z(n1928) );
  IVSVTX4 U1850 ( .A(n514), .Z(n3147) );
  CTIVSVTX2 U1851 ( .A(n989), .Z(n3601) );
  CTIVSVTX2 U1852 ( .A(n3183), .Z(n3187) );
  ND2SVTX2 U1853 ( .A(n3114), .B(n4134), .Z(n887) );
  IVSVTX10 U1854 ( .A(n2424), .Z(n4073) );
  AO1ASVTX6 U1855 ( .A(n3332), .B(n4151), .C(n3123), .D(n1575), .Z(n4153) );
  ND2SVTX4 U1856 ( .A(n4099), .B(n3142), .Z(n4139) );
  CTIVSVTX4 U1857 ( .A(n480), .Z(n2276) );
  IVSVTX4 U1858 ( .A(n3739), .Z(n526) );
  ND3SVTX4 U1859 ( .A(n1132), .B(n3620), .C(n880), .Z(n1129) );
  NR2SVTX4 U1860 ( .A(n3797), .B(n583), .Z(n1338) );
  ND2SVTX4 U1861 ( .A(n1966), .B(n3984), .Z(n1850) );
  IVSVTX8 U1862 ( .A(n697), .Z(n530) );
  IVSVTX8 U1863 ( .A(n4179), .Z(n509) );
  NR2SVTX2 U1864 ( .A(n474), .B(n1878), .Z(n1649) );
  ND2SVTX2 U1865 ( .A(n3711), .B(n1428), .Z(n1470) );
  IVSVTX4 U1866 ( .A(n2936), .Z(n4070) );
  CTIVSVTX4 U1867 ( .A(n1869), .Z(n3937) );
  ND3SVTX4 U1868 ( .A(n2442), .B(n531), .C(n3203), .Z(n1486) );
  IVSVTX4 U1869 ( .A(n1878), .Z(n3739) );
  ND3ABSVTX4 U1870 ( .A(n3878), .B(n3874), .C(n876), .Z(n3877) );
  NR2ASVTX2 U1871 ( .A(n3693), .B(n3627), .Z(n3630) );
  B_ND2SVTX2 U1872 ( .A(n4163), .B(n4150), .Z(n4108) );
  AO6SVTX4 U1873 ( .A(n3982), .B(n2913), .C(n1220), .Z(n3237) );
  IVSVTX2 U1874 ( .A(n3245), .Z(n1922) );
  IVSVTX2 U1875 ( .A(n1176), .Z(n3989) );
  CTIVSVTX4 U1876 ( .A(n3498), .Z(n3499) );
  IVSVTX2 U1877 ( .A(n660), .Z(n1877) );
  CTIVSVTX2 U1878 ( .A(n2866), .Z(n2926) );
  IVSVTX4 U1879 ( .A(n1719), .Z(n3105) );
  AO7ABSVTX6 U1880 ( .A(n507), .B(n2781), .C(n2780), .Z(n2938) );
  CTIVSVTX2 U1881 ( .A(n1839), .Z(n1970) );
  IVSVTX4 U1882 ( .A(n3212), .Z(n780) );
  AO7ABSVTX6 U1883 ( .A(n610), .B(n507), .C(n2770), .Z(n1745) );
  ND3SVTX6 U1884 ( .A(n2830), .B(n1325), .C(n1326), .Z(n3719) );
  ND2SVTX2 U1885 ( .A(n3980), .B(n1177), .Z(n1176) );
  ND2SVTX4 U1886 ( .A(n2050), .B(n1840), .Z(n3623) );
  IVSVTX6 U1887 ( .A(n2805), .Z(n2770) );
  CTIVSVTX2 U1888 ( .A(n2399), .Z(n1689) );
  B_ND2SVTX2 U1889 ( .A(n3852), .B(n3853), .Z(n3858) );
  IVSVTX2 U1890 ( .A(n3432), .Z(n2035) );
  IVSVTX2 U1891 ( .A(n1615), .Z(n3520) );
  IVSVTX4 U1892 ( .A(n3706), .Z(n595) );
  AN2SVTX4 U1893 ( .A(n2328), .B(n3029), .Z(n3123) );
  F_IVSVTX1 U1894 ( .A(n2454), .Z(n1608) );
  ND2SVTX2 U1895 ( .A(n2808), .B(n610), .Z(n1416) );
  IVSVTX2 U1896 ( .A(n2742), .Z(n1671) );
  ND2SVTX8 U1897 ( .A(n2052), .B(n3621), .Z(n2050) );
  IVSVTX2 U1898 ( .A(n3121), .Z(n3125) );
  NR2SVTX4 U1899 ( .A(n2052), .B(n3621), .Z(n1326) );
  ND2SVTX4 U1900 ( .A(n3054), .B(n3053), .Z(n4035) );
  CTIVSVTX4 U1901 ( .A(n2897), .Z(n2909) );
  AN2SVTX6 U1902 ( .A(n3006), .B(n3005), .Z(n1079) );
  ND2SVTX6 U1903 ( .A(n604), .B(n1080), .Z(n3973) );
  IVSVTX2 U1904 ( .A(n3099), .Z(n3049) );
  ND2ASVTX6 U1905 ( .A(n2891), .B(n613), .Z(n3662) );
  AO7ABSVTX6 U1906 ( .A(n541), .B(n1006), .C(n1355), .Z(n2815) );
  NR2ASVTX2 U1907 ( .A(n2347), .B(n3639), .Z(n3604) );
  ND2SVTX2 U1908 ( .A(n1333), .B(n1331), .Z(n2808) );
  CTIVSVTX2 U1909 ( .A(n3935), .Z(n2301) );
  ND2SVTX4 U1910 ( .A(n2918), .B(n2917), .Z(n3853) );
  ENSVTX6 U1911 ( .A(n1828), .B(n2844), .Z(n3442) );
  IVSVTX4 U1912 ( .A(n948), .Z(n608) );
  ND2SVTX2 U1913 ( .A(n444), .B(n1332), .Z(n1331) );
  ND2SVTX2 U1914 ( .A(n1226), .B(n1224), .Z(n3010) );
  IVSVTX4 U1915 ( .A(n3287), .Z(n517) );
  AO7SVTX4 U1916 ( .A(n3495), .B(n3284), .C(n3493), .Z(n3434) );
  ND2SVTX4 U1917 ( .A(n1814), .B(n1813), .Z(n2891) );
  ND2SVTX4 U1918 ( .A(n808), .B(n687), .Z(n816) );
  B_ND2SVTX1 U1919 ( .A(n3478), .B(n3477), .Z(n3480) );
  CTIVSVTX2 U1920 ( .A(n3494), .Z(n3284) );
  ND2SVTX6 U1921 ( .A(n1569), .B(n1853), .Z(n1536) );
  IVSVTX10 U1922 ( .A(n1389), .Z(n542) );
  IVSVTX8 U1923 ( .A(n1480), .Z(n1481) );
  ND2SVTX6 U1924 ( .A(n1000), .B(n1048), .Z(n1389) );
  ND2SVTX6 U1925 ( .A(n2674), .B(n2675), .Z(n683) );
  ND2SVTX6 U1926 ( .A(n549), .B(n2610), .Z(n2619) );
  NR3ABSVTX6 U1927 ( .A(n2132), .B(n1096), .C(n1095), .Z(n2613) );
  ND2ASVTX4 U1928 ( .A(n2671), .B(n1904), .Z(n2537) );
  IVSVTX2 U1929 ( .A(n2622), .Z(n1773) );
  ND3ASVTX6 U1930 ( .A(n555), .B(n1904), .C(n2231), .Z(n2563) );
  IVSVTX4 U1931 ( .A(n2364), .Z(n1805) );
  IVSVTX8 U1932 ( .A(n2571), .Z(n513) );
  IVSVTX4 U1933 ( .A(num_i[10]), .Z(n553) );
  OR2SVTX4 U1934 ( .A(n4188), .B(n1659), .Z(n4186) );
  B_ND2SVTX2 U1935 ( .A(n4220), .B(n4219), .Z(n4223) );
  IVSVTX2 U1936 ( .A(n4277), .Z(n1465) );
  NR2SVTX4 U1937 ( .A(n4111), .B(n1925), .Z(n4112) );
  B_ND2SVTX2 U1938 ( .A(n4183), .B(n4182), .Z(n2304) );
  F_AN2SVTX2 U1939 ( .A(n4213), .B(n2368), .Z(n2447) );
  ND3SVTX4 U1940 ( .A(n1926), .B(n1350), .C(n1930), .Z(n1925) );
  ND2SVTX2 U1941 ( .A(n2122), .B(n2121), .Z(n2042) );
  B_ND2SVTX2 U1942 ( .A(n4244), .B(n4235), .Z(n4246) );
  NR3ABSVTX4 U1943 ( .A(n1012), .B(n2445), .C(n1010), .Z(n1795) );
  IVSVTX2 U1944 ( .A(n764), .Z(n1456) );
  ND3ABSVTX4 U1945 ( .A(n3977), .B(n3974), .C(n557), .Z(n2028) );
  ND3ASVTX6 U1946 ( .A(n4048), .B(n1012), .C(n1673), .Z(n1011) );
  NR2SVTX6 U1947 ( .A(n566), .B(n954), .Z(n4234) );
  AO7SVTX2 U1948 ( .A(n3210), .B(n3209), .C(n733), .Z(n2123) );
  F_AN2SVTX2 U1949 ( .A(n2767), .B(n2766), .Z(n2768) );
  ND3SVTX4 U1950 ( .A(n3946), .B(n3947), .C(n2359), .Z(n1193) );
  AO6SVTX2 U1951 ( .A(n838), .B(n2451), .C(n837), .Z(n1918) );
  AO7SVTX2 U1952 ( .A(n3601), .B(n3600), .C(n733), .Z(n3602) );
  CTIVSVTX10 U1953 ( .A(n3117), .Z(n3260) );
  IVSVTX4 U1954 ( .A(n739), .Z(n4160) );
  AO7ASVTX4 U1955 ( .A(n753), .B(n1525), .C(n3989), .Z(n3990) );
  ND3SVTX2 U1956 ( .A(n733), .B(n2031), .C(n2030), .Z(n2029) );
  OR2SVTX4 U1957 ( .A(n526), .B(n3368), .Z(n2426) );
  ND2SVTX2 U1958 ( .A(n1789), .B(n2103), .Z(n766) );
  CTIVSVTX2 U1959 ( .A(n3230), .Z(n3231) );
  IVSVTX2 U1960 ( .A(n3430), .Z(n1100) );
  ND3SVTX4 U1961 ( .A(n3135), .B(n865), .C(n3134), .Z(n2086) );
  IVSVTX4 U1962 ( .A(n3983), .Z(n569) );
  AO2SVTX4 U1963 ( .A(n3605), .B(n530), .C(n823), .D(n441), .Z(n3701) );
  ND3SVTX2 U1964 ( .A(n468), .B(n1471), .C(n1470), .Z(n3708) );
  CTIVSVTX2 U1965 ( .A(n3156), .Z(n3157) );
  ND2ASVTX4 U1966 ( .A(n1627), .B(n530), .Z(n1950) );
  NR3ABSVTX4 U1967 ( .A(n3489), .B(n3429), .C(n3490), .Z(n3430) );
  ND3SVTX4 U1968 ( .A(n4150), .B(n740), .C(n4151), .Z(n739) );
  IVSVTX2 U1969 ( .A(n3402), .Z(n3403) );
  NR2ASVTX4 U1970 ( .A(n530), .B(n2315), .Z(n2079) );
  ND2SVTX2 U1971 ( .A(n3977), .B(n3978), .Z(n2030) );
  CTIVSVTX2 U1972 ( .A(n3978), .Z(n3979) );
  AO2SVTX2 U1973 ( .A(n3697), .B(n3696), .C(n2354), .D(n3695), .Z(n1750) );
  B_ND2SVTX2 U1974 ( .A(n3976), .B(n3975), .Z(n2031) );
  IVSVTX4 U1975 ( .A(n830), .Z(n831) );
  CTIVSVTX2 U1976 ( .A(n3239), .Z(n3229) );
  B_ND2SVTX2 U1977 ( .A(n3148), .B(n4121), .Z(n3156) );
  AO6SVTX2 U1978 ( .A(n3031), .B(n3030), .C(n3124), .Z(n1575) );
  CTBUFSVTX12 U1979 ( .A(n648), .Z(n1422) );
  B_ND2SVTX2 U1980 ( .A(n3707), .B(n3709), .Z(n1471) );
  B_ND2SVTX2 U1981 ( .A(n3679), .B(n3678), .Z(n1386) );
  CTIVSVTX2 U1982 ( .A(n3141), .Z(n1283) );
  IVSVTX6 U1983 ( .A(n3951), .Z(n533) );
  NR2SVTX6 U1984 ( .A(n3421), .B(n1077), .Z(n3427) );
  AO7ABSVTX2 U1985 ( .A(n3126), .B(n3121), .C(n1922), .Z(n3031) );
  NR3ABSVTX6 U1986 ( .A(n3420), .B(n3973), .C(n3977), .Z(n991) );
  AO6SVTX4 U1987 ( .A(n1994), .B(n4009), .C(n3292), .Z(n3344) );
  IVSVTX4 U1988 ( .A(n3325), .Z(n531) );
  IVSVTX2 U1989 ( .A(n3545), .Z(n3540) );
  ND4ABSVTX6 U1990 ( .A(n510), .B(n1148), .C(n3663), .D(n1040), .Z(n2242) );
  IVSVTX4 U1991 ( .A(n1824), .Z(n576) );
  IVSVTX2 U1992 ( .A(n536), .Z(n2224) );
  IVSVTX4 U1993 ( .A(n1513), .Z(n1146) );
  ND2SVTX4 U1994 ( .A(n2979), .B(n2980), .Z(n2379) );
  ND2ASVTX6 U1995 ( .A(n1751), .B(n1286), .Z(n4055) );
  IVSVTX2 U1996 ( .A(n3684), .Z(n3685) );
  AO17SVTX4 U1997 ( .A(n1053), .B(n2959), .C(n3372), .D(n3267), .Z(n3325) );
  CTIVSVTX2 U1998 ( .A(n3419), .Z(n2326) );
  B_ND2SVTX2 U1999 ( .A(n3034), .B(n3033), .Z(n4152) );
  F_ND2ASVTX2 U2000 ( .A(n3533), .B(n3532), .Z(n3535) );
  IVSVTX2 U2001 ( .A(n2826), .Z(n2827) );
  NR2ASVTX4 U2002 ( .A(n3691), .B(n2997), .Z(n3597) );
  IVSVTX2 U2003 ( .A(n3612), .Z(n924) );
  CTIVSVTX2 U2004 ( .A(n3889), .Z(n3829) );
  CTBUFSVTX4 U2005 ( .A(n3590), .Z(n1617) );
  CTAN2BSVTX4 U2006 ( .A(n3365), .B(n3048), .Z(n3368) );
  ND2SVTX4 U2007 ( .A(n2904), .B(n2903), .Z(n2358) );
  ND2ASVTX6 U2008 ( .A(n3504), .B(n1606), .Z(n3524) );
  IVSVTX4 U2009 ( .A(n2917), .Z(n2904) );
  B_ND2SVTX2 U2010 ( .A(n1790), .B(n606), .Z(n4120) );
  ND2SVTX4 U2011 ( .A(n2906), .B(n1595), .Z(n2910) );
  IVSVTX4 U2012 ( .A(n1058), .Z(n1059) );
  ND2ASVTX4 U2013 ( .A(n543), .B(n1523), .Z(n3288) );
  IVSVTX2 U2014 ( .A(n2798), .Z(n1581) );
  IVSVTX6 U2015 ( .A(n2865), .Z(n2945) );
  ND2SVTX2 U2016 ( .A(n1961), .B(n3668), .Z(n1960) );
  NR2ASVTX2 U2017 ( .A(n3516), .B(n3515), .Z(n3517) );
  NR2SVTX2 U2018 ( .A(n4005), .B(n4004), .Z(n4017) );
  NR2ASVTX6 U2019 ( .A(n3079), .B(n3075), .Z(n1623) );
  IVSVTX2 U2020 ( .A(n3672), .Z(n1961) );
  IVSVTX8 U2021 ( .A(n2128), .Z(n518) );
  IVSVTX6 U2022 ( .A(n3282), .Z(n1881) );
  IVSVTX8 U2023 ( .A(n628), .Z(n643) );
  F_IVSVTX1 U2024 ( .A(n508), .Z(n1033) );
  IVSVTX4 U2025 ( .A(n681), .Z(n1534) );
  IVSVTX12 U2026 ( .A(n1770), .Z(n519) );
  AO7SVTX4 U2027 ( .A(n634), .B(n2332), .C(n968), .Z(n1056) );
  ND2SVTX6 U2028 ( .A(n1034), .B(n1039), .Z(n2549) );
  IVSVTX2 U2029 ( .A(n2415), .Z(n1677) );
  AN2SVTX4 U2030 ( .A(n552), .B(n2672), .Z(n2627) );
  ND3ABSVTX4 U2031 ( .A(n656), .B(n657), .C(n512), .Z(n2626) );
  NR2ASVTX4 U2032 ( .A(n1755), .B(rslt_o[31]), .Z(n2689) );
  IVSVTX2 U2033 ( .A(n1805), .Z(n657) );
  IVSVTX2 U2034 ( .A(n2635), .Z(n2622) );
  IVSVTX2 U2035 ( .A(n2369), .Z(n913) );
  IVSVTX4 U2036 ( .A(n2696), .Z(n550) );
  ND2SVTX4 U2037 ( .A(n2492), .B(n2499), .Z(n2495) );
  CTIVSVTX2 U2038 ( .A(n2644), .Z(n1723) );
  CTIVSVTX2 U2039 ( .A(n2624), .Z(n2517) );
  CTIVSVTX2 U2040 ( .A(n554), .Z(n2013) );
  CTBUFSVTX4 U2041 ( .A(num_i[7]), .Z(n2638) );
  CTIVSVTX4 U2042 ( .A(n4205), .Z(n4194) );
  ENSVTX4 U2043 ( .A(n4243), .B(n4301), .Z(rslt_o[9]) );
  B_ND2SVTX2 U2044 ( .A(n3110), .B(n3109), .Z(n4090) );
  IVSVTX2 U2045 ( .A(n4292), .Z(n1626) );
  EOSVTX4 U2046 ( .A(n4246), .B(n4245), .Z(rslt_o[6]) );
  ND2SVTX6 U2047 ( .A(n1009), .B(n2357), .Z(n4219) );
  ENSVTX4 U2048 ( .A(n4256), .B(n4255), .Z(rslt_o[4]) );
  B_ND2SVTX2 U2049 ( .A(n4277), .B(n412), .Z(n4280) );
  ENSVTX4 U2050 ( .A(n1722), .B(n4259), .Z(rslt_o[3]) );
  IVSVTX4 U2051 ( .A(n1014), .Z(n2357) );
  NR2SVTX2 U2052 ( .A(n2304), .B(n2302), .Z(n4184) );
  ND2SVTX4 U2053 ( .A(n2040), .B(n2042), .Z(n2039) );
  ND2SVTX4 U2054 ( .A(n1946), .B(n4229), .Z(n3687) );
  B_ND2SVTX1 U2055 ( .A(n4229), .B(n4230), .Z(n4233) );
  IVSVTX6 U2056 ( .A(n2368), .Z(n1914) );
  ND3ABSVTX4 U2057 ( .A(n1983), .B(n3383), .C(n4095), .Z(n4114) );
  ND3ABSVTX6 U2058 ( .A(n1519), .B(n490), .C(n1746), .Z(n4113) );
  ND2SVTX4 U2059 ( .A(n3854), .B(n1403), .Z(n4288) );
  AO1ABSVTX4 U2060 ( .A(n597), .B(n4109), .C(n4180), .D(n1752), .Z(n4111) );
  IVSVTX2 U2061 ( .A(n3159), .Z(n1356) );
  B_ND2SVTX2 U2062 ( .A(n4170), .B(n4169), .Z(n4185) );
  ND2ASVTX4 U2063 ( .A(n2029), .B(n2028), .Z(n3994) );
  NR3ABSVTX4 U2064 ( .A(n3347), .B(n1596), .C(n2277), .Z(n1414) );
  ND3SVTX6 U2065 ( .A(n2411), .B(n3602), .C(n3617), .Z(n4229) );
  IVSVTX2 U2066 ( .A(n2123), .Z(n2122) );
  CTIVSVTX2 U2067 ( .A(n2356), .Z(n4173) );
  IVSVTX2 U2068 ( .A(n2165), .Z(n1752) );
  ND3SVTX4 U2069 ( .A(n1415), .B(n1412), .C(n2274), .Z(n1411) );
  ND4ABSVTX4 U2070 ( .A(n3231), .B(n3232), .C(n2091), .D(n1172), .Z(n2090) );
  ND4ASVTX4 U2071 ( .A(n1614), .B(n3253), .C(n3332), .D(n3252), .Z(n3255) );
  IVSVTX6 U2072 ( .A(n960), .Z(n557) );
  CTIVSVTX4 U2073 ( .A(n2234), .Z(n1843) );
  ND3SVTX4 U2074 ( .A(n2114), .B(n1596), .C(n1190), .Z(n1189) );
  ND2SVTX4 U2075 ( .A(n1632), .B(n2310), .Z(n1182) );
  NR3ABSVTX4 U2076 ( .A(n3427), .B(n3425), .C(n960), .Z(n2188) );
  ND2SVTX4 U2077 ( .A(n1181), .B(n1193), .Z(n1180) );
  AO7SVTX4 U2078 ( .A(n1574), .B(n1573), .C(n1422), .Z(n1930) );
  ND3ABSVTX4 U2079 ( .A(n3427), .B(n3426), .C(n960), .Z(n2187) );
  NR2SVTX4 U2080 ( .A(n3979), .B(n557), .Z(n3993) );
  NR2SVTX4 U2081 ( .A(n1779), .B(n4126), .Z(n1778) );
  ND4ABSVTX6 U2082 ( .A(n3116), .B(n2113), .C(n4091), .D(n3146), .Z(n1468) );
  ND2SVTX4 U2083 ( .A(n2410), .B(n2124), .Z(n2047) );
  AO7ABSVTX2 U2084 ( .A(n4046), .B(n4045), .C(n4044), .Z(n4047) );
  IVSVTX4 U2085 ( .A(n868), .Z(n867) );
  NR2ASVTX4 U2086 ( .A(n2201), .B(n560), .Z(n1713) );
  B_ND2SVTX2 U2087 ( .A(n506), .B(n4126), .Z(n4129) );
  NR4ABSVTX6 U2088 ( .A(n3971), .B(n1196), .C(n1194), .D(n1185), .Z(n1181) );
  IVSVTX4 U2089 ( .A(n1533), .Z(n1876) );
  ND3SVTX4 U2090 ( .A(n2276), .B(n838), .C(n1405), .Z(n1404) );
  ND3ABSVTX6 U2091 ( .A(n3849), .B(n1754), .C(n1753), .Z(n3850) );
  NR2SVTX4 U2092 ( .A(n3801), .B(n3800), .Z(n3805) );
  IVSVTX4 U2093 ( .A(n1485), .Z(n788) );
  ND2ASVTX4 U2094 ( .A(n1635), .B(n3376), .Z(n3375) );
  AO7SVTX4 U2095 ( .A(n3419), .B(n1900), .C(n1899), .Z(n1898) );
  NR3ASVTX6 U2096 ( .A(n568), .B(n2426), .C(n562), .Z(n1920) );
  ND3ABSVTX4 U2097 ( .A(n1635), .B(n3377), .C(n3376), .Z(n3378) );
  IVSVTX2 U2098 ( .A(n1706), .Z(n3904) );
  ND3SVTX6 U2099 ( .A(n2229), .B(n3902), .C(n2340), .Z(n868) );
  AO7NSVTX2 U2100 ( .A(n3716), .B(n2413), .C(n566), .Z(n2383) );
  NR2SVTX4 U2101 ( .A(n1214), .B(n1211), .Z(n1104) );
  CTIVSVTX2 U2102 ( .A(n2828), .Z(n2943) );
  AO7SVTX2 U2103 ( .A(n2233), .B(n1750), .C(n2293), .Z(n3698) );
  AO7SVTX4 U2104 ( .A(n3330), .B(n3328), .C(n733), .Z(n1485) );
  IVSVTX10 U2105 ( .A(n769), .Z(n3179) );
  AO1SVTX4 U2106 ( .A(n3732), .B(n3731), .C(n3729), .D(n3730), .Z(n3733) );
  IVSVTX2 U2107 ( .A(n766), .Z(n3389) );
  ND3SVTX4 U2108 ( .A(n1213), .B(n3482), .C(n1212), .Z(n1211) );
  IVSVTX8 U2109 ( .A(n4075), .Z(n3164) );
  IVSVTX8 U2110 ( .A(n1367), .Z(n1246) );
  AO7SVTX4 U2111 ( .A(n4101), .B(n1243), .C(n572), .Z(n1161) );
  B_ND2SVTX2 U2112 ( .A(n3184), .B(n3187), .Z(n3197) );
  CTBUFSVTX4 U2113 ( .A(n3905), .Z(n1706) );
  AO4SVTX4 U2114 ( .A(n3999), .B(n3383), .C(n3383), .D(n1173), .Z(n4003) );
  NR2SVTX6 U2115 ( .A(n733), .B(n514), .Z(n2394) );
  IVSVTX2 U2116 ( .A(n3699), .Z(n1818) );
  ND3ABSVTX4 U2117 ( .A(n1690), .B(n2291), .C(n990), .Z(n3699) );
  NR2ASVTX4 U2118 ( .A(n585), .B(n3732), .Z(n3730) );
  IVSVTX2 U2119 ( .A(n3714), .Z(n1820) );
  ND2ASVTX6 U2120 ( .A(n2292), .B(n4050), .Z(n1866) );
  ND3ABSVTX4 U2121 ( .A(n1591), .B(n4092), .C(n2418), .Z(n2055) );
  ND2SVTX4 U2122 ( .A(n1951), .B(n1950), .Z(n1949) );
  NR3SVTX4 U2123 ( .A(n515), .B(n4073), .C(n1376), .Z(n1375) );
  AO1ASVTX4 U2124 ( .A(n2050), .B(n3903), .C(n4073), .D(n1969), .Z(n1968) );
  ND3SVTX4 U2125 ( .A(n3769), .B(n1883), .C(n3771), .Z(n3778) );
  AO3SVTX4 U2126 ( .A(n1838), .B(n3951), .C(n1422), .D(n4036), .Z(n1880) );
  NR3SVTX4 U2127 ( .A(n4073), .B(n3842), .C(n3847), .Z(n3843) );
  AO4SVTX4 U2128 ( .A(n3686), .B(n455), .C(n2380), .D(n2351), .Z(n2254) );
  AO6ABSVTX6 U2129 ( .A(n1507), .B(n576), .C(n866), .Z(n3470) );
  ND4SVTX4 U2130 ( .A(n1218), .B(n648), .C(n1217), .D(n1216), .Z(n1212) );
  ND2SVTX4 U2131 ( .A(n1487), .B(n1486), .Z(n3328) );
  F_ENSVTX2 U2132 ( .A(n3388), .B(n3387), .Z(n2236) );
  IVSVTX8 U2133 ( .A(n907), .Z(n1740) );
  CTIVSVTX2 U2134 ( .A(n3178), .Z(n3181) );
  ND2ASVTX4 U2135 ( .A(n1288), .B(n1289), .Z(n3230) );
  IVSVTX12 U2136 ( .A(n4066), .Z(n524) );
  CTIVSVTX4 U2137 ( .A(n2056), .Z(n2418) );
  ND3SVTX4 U2138 ( .A(n2064), .B(n3484), .C(n745), .Z(n848) );
  ND2SVTX2 U2139 ( .A(n402), .B(n441), .Z(n4019) );
  IVSVTX2 U2140 ( .A(n1497), .Z(n1490) );
  IVSVTX4 U2141 ( .A(n1132), .Z(n1131) );
  NR2SVTX2 U2142 ( .A(n1448), .B(n3713), .Z(n3714) );
  ND2SVTX4 U2143 ( .A(n1495), .B(n1494), .Z(n1493) );
  IVSVTX4 U2144 ( .A(n1635), .Z(n567) );
  AO7SVTX4 U2145 ( .A(n3823), .B(n3822), .C(n648), .Z(n1424) );
  B_ND2SVTX2 U2146 ( .A(n2424), .B(n457), .Z(n2756) );
  IVSVTX2 U2147 ( .A(n3692), .Z(n990) );
  IVSVTX2 U2148 ( .A(n3696), .Z(n3692) );
  AO7SVTX2 U2149 ( .A(n3875), .B(n3874), .C(n3878), .Z(n3876) );
  IVSVTX2 U2150 ( .A(n4117), .Z(n1725) );
  IVSVTX8 U2151 ( .A(n2292), .Z(n2291) );
  IVSVTX8 U2152 ( .A(n3162), .Z(n528) );
  IVSVTX8 U2153 ( .A(n3211), .Z(n570) );
  AO7SVTX4 U2154 ( .A(n611), .B(n3112), .C(n2393), .Z(n1549) );
  B_ND2SVTX2 U2155 ( .A(n582), .B(n3239), .Z(n3225) );
  NR2ASVTX6 U2156 ( .A(n1498), .B(n2058), .Z(n1497) );
  AO7SVTX4 U2157 ( .A(n584), .B(n1192), .C(n3722), .Z(n3962) );
  NR2ASVTX4 U2158 ( .A(n2397), .B(n3753), .Z(n3754) );
  IVSVTX4 U2159 ( .A(n3206), .Z(n3012) );
  IVSVTX2 U2160 ( .A(n3336), .Z(n2027) );
  NR3SVTX4 U2161 ( .A(n906), .B(n3831), .C(n697), .Z(n3833) );
  NR2SVTX6 U2162 ( .A(n3072), .B(n3071), .Z(n3814) );
  CTIVSVTX2 U2163 ( .A(n515), .Z(n3659) );
  AO7SVTX4 U2164 ( .A(n2224), .B(n3998), .C(n1409), .Z(n957) );
  CTIVSVTX2 U2165 ( .A(n3657), .Z(n1376) );
  NR3ABSVTX6 U2166 ( .A(n3021), .B(n2119), .C(n1877), .Z(n1878) );
  IVSVTX8 U2167 ( .A(n1016), .Z(n3795) );
  NR2SVTX6 U2168 ( .A(n3811), .B(n3087), .Z(n2205) );
  ND3ASVTX6 U2169 ( .A(n3745), .B(n4014), .C(n1994), .Z(n3343) );
  AO6SVTX2 U2170 ( .A(n3611), .B(n924), .C(n922), .Z(n921) );
  AO6SVTX6 U2171 ( .A(n3586), .B(n3587), .C(n3585), .Z(n3629) );
  IVSVTX4 U2172 ( .A(n3690), .Z(n830) );
  NR2SVTX2 U2173 ( .A(n3989), .B(n3982), .Z(n1524) );
  AO7SVTX4 U2174 ( .A(n590), .B(n481), .C(n1177), .Z(n3417) );
  ND2SVTX6 U2175 ( .A(n3367), .B(n1364), .Z(n4057) );
  IVSVTX4 U2176 ( .A(n4039), .Z(n1302) );
  IVSVTX2 U2177 ( .A(n3678), .Z(n3669) );
  AO7ASVTX6 U2178 ( .A(n803), .B(n805), .C(n3084), .Z(n806) );
  ND2SVTX4 U2179 ( .A(n1066), .B(n2152), .Z(n1065) );
  IVSVTX4 U2180 ( .A(n1856), .Z(n1387) );
  NR2SVTX4 U2181 ( .A(n3087), .B(n3064), .Z(n3171) );
  IVSVTX4 U2182 ( .A(n3770), .Z(n3771) );
  ND2ASVTX4 U2183 ( .A(n3870), .B(n3879), .Z(n3824) );
  IVSVTX4 U2184 ( .A(n3223), .Z(n581) );
  ND3SVTX6 U2185 ( .A(n3738), .B(n3787), .C(n3933), .Z(n4039) );
  NR2ASVTX4 U2186 ( .A(n1839), .B(n3903), .Z(n1969) );
  IVSVTX4 U2187 ( .A(n3462), .Z(n577) );
  AO7SVTX4 U2188 ( .A(n1324), .B(n1840), .C(n1499), .Z(n3842) );
  ND2ASVTX4 U2189 ( .A(n755), .B(n3888), .Z(n926) );
  ND2ASVTX6 U2190 ( .A(n3122), .B(n2946), .Z(n4121) );
  AO7SVTX6 U2191 ( .A(n1808), .B(n3489), .C(n3428), .Z(n3585) );
  ND2SVTX4 U2192 ( .A(n1943), .B(n1944), .Z(n1942) );
  MUX21NSVTX2 U2193 ( .A(n3489), .B(n1617), .S(n3429), .Z(n3431) );
  IVSVTX4 U2194 ( .A(n3374), .Z(n3324) );
  AO7SVTX4 U2195 ( .A(n610), .B(n3310), .C(n1719), .Z(n2437) );
  NR2ASVTX4 U2196 ( .A(n3489), .B(n588), .Z(n3491) );
  CTIVSVTX2 U2197 ( .A(n3276), .Z(n3277) );
  ND2SVTX6 U2198 ( .A(n2895), .B(n3772), .Z(n3690) );
  ND2SVTX6 U2199 ( .A(n3840), .B(n1017), .Z(n1016) );
  CTIVSVTX4 U2200 ( .A(n3170), .Z(n534) );
  IVSVTX4 U2201 ( .A(n3745), .Z(n3939) );
  IVSVTX4 U2202 ( .A(n2020), .Z(n1934) );
  CTIVSVTX4 U2203 ( .A(n3969), .Z(n535) );
  ND2SVTX4 U2204 ( .A(n3086), .B(n1915), .Z(n1944) );
  B_ND2SVTX2 U2205 ( .A(n615), .B(n4135), .Z(n4172) );
  CTIVSVTX2 U2206 ( .A(n415), .Z(n4034) );
  IVSVTX2 U2207 ( .A(n3656), .Z(n3655) );
  NR2SVTX2 U2208 ( .A(n3684), .B(n3597), .Z(n3598) );
  ND3SVTX4 U2209 ( .A(n3846), .B(n644), .C(n511), .Z(n1663) );
  ND2SVTX2 U2210 ( .A(n3612), .B(n3610), .Z(n923) );
  IVSVTX4 U2211 ( .A(n1617), .Z(n588) );
  ND2ASVTX4 U2212 ( .A(n2341), .B(n2343), .Z(n2716) );
  ND2SVTX4 U2213 ( .A(n3457), .B(n1551), .Z(n3462) );
  NR2SVTX6 U2214 ( .A(n2925), .B(n2924), .Z(n3223) );
  ENSVTX4 U2215 ( .A(n2776), .B(n1577), .Z(n2946) );
  IVSVTX4 U2216 ( .A(n3857), .Z(n801) );
  IVSVTX4 U2217 ( .A(n2216), .Z(n1286) );
  CTIVSVTX2 U2218 ( .A(n1257), .Z(n1256) );
  IVSVTX2 U2219 ( .A(n3175), .Z(n3127) );
  CTIVSVTX4 U2220 ( .A(n1079), .Z(n3955) );
  B_ND2SVTX2 U2221 ( .A(n3412), .B(n3411), .Z(n3419) );
  ND2ASVTX6 U2222 ( .A(n599), .B(n2089), .Z(n1177) );
  ND2ASVTX4 U2223 ( .A(n2776), .B(n1671), .Z(n2744) );
  IVSVTX4 U2224 ( .A(n1004), .Z(n536) );
  NR2ASVTX4 U2225 ( .A(n3893), .B(n3898), .Z(n3895) );
  IVSVTX2 U2226 ( .A(n3289), .Z(n3291) );
  AO7SVTX6 U2227 ( .A(n2719), .B(n2708), .C(n2776), .Z(n2715) );
  IVSVTX8 U2228 ( .A(n821), .Z(n3589) );
  NR2SVTX6 U2229 ( .A(n3080), .B(n3501), .Z(n1915) );
  AO7SVTX2 U2230 ( .A(n4006), .B(n2158), .C(n2156), .Z(n3292) );
  CTIVSVTX2 U2231 ( .A(n3524), .Z(n3523) );
  IVSVTX2 U2232 ( .A(n3007), .Z(n3009) );
  CTBUFSVTX4 U2233 ( .A(n3552), .Z(n799) );
  NR2SVTX6 U2234 ( .A(n2996), .B(n603), .Z(n821) );
  AO7SVTX4 U2235 ( .A(n2199), .B(n3270), .C(n1791), .Z(n2977) );
  NR2ASVTX4 U2236 ( .A(n3111), .B(n3121), .Z(n1638) );
  ND2ASVTX4 U2237 ( .A(n3111), .B(n3121), .Z(n3175) );
  IVSVTX4 U2238 ( .A(n2910), .Z(n599) );
  IVSVTX4 U2239 ( .A(n3583), .Z(n2997) );
  AO7ABSVTX6 U2240 ( .A(n2868), .B(n1482), .C(n2215), .Z(n2781) );
  IVSVTX2 U2241 ( .A(n3288), .Z(n3533) );
  ND2SVTX4 U2242 ( .A(n1837), .B(n3058), .Z(n3095) );
  NR2ASVTX6 U2243 ( .A(n2798), .B(n2800), .Z(n2935) );
  IVSVTX2 U2244 ( .A(n3554), .Z(n3510) );
  AO7SVTX4 U2245 ( .A(n2807), .B(n1571), .C(n2945), .Z(n1578) );
  AO7ABSVTX4 U2246 ( .A(n606), .B(n3270), .C(n1294), .Z(n3040) );
  ND2ASVTX6 U2247 ( .A(n506), .B(n2787), .Z(n2777) );
  CTIVSVTX2 U2248 ( .A(n2927), .Z(n2867) );
  ND2SVTX6 U2249 ( .A(n2821), .B(n2823), .Z(n2830) );
  ND2SVTX6 U2250 ( .A(n607), .B(n2876), .Z(n3703) );
  B_ND2SVTX2 U2251 ( .A(n3285), .B(n3287), .Z(n2747) );
  ND2SVTX6 U2252 ( .A(n1921), .B(n3958), .Z(n3880) );
  ND2SVTX6 U2253 ( .A(n2710), .B(n2709), .Z(n2711) );
  AO4SVTX6 U2254 ( .A(n2785), .B(n606), .C(n617), .D(n1790), .Z(n2790) );
  AN3SVTX6 U2255 ( .A(n2348), .B(n608), .C(n2309), .Z(n2087) );
  B_ND2SVTX2 U2256 ( .A(n871), .B(n3505), .Z(n2759) );
  OR2SVTX4 U2257 ( .A(n2745), .B(n3451), .Z(n2746) );
  ND2ASVTX6 U2258 ( .A(n3459), .B(n3083), .Z(n3471) );
  ND2SVTX6 U2259 ( .A(n2460), .B(n2404), .Z(n3959) );
  IVSVTX2 U2260 ( .A(n2743), .Z(n1088) );
  IVSVTX4 U2261 ( .A(n3091), .Z(n3061) );
  CTIVSVTX4 U2262 ( .A(n2988), .Z(n603) );
  IVSVTX2 U2263 ( .A(n2717), .Z(n2718) );
  ND2SVTX6 U2264 ( .A(n3063), .B(n3062), .Z(n3607) );
  F_ENSVTX2 U2265 ( .A(n1547), .B(n2344), .Z(n2955) );
  ND2SVTX6 U2266 ( .A(n2719), .B(n759), .Z(n2288) );
  AO5NSVTX4 U2267 ( .A(n652), .B(n2807), .C(n621), .Z(n1751) );
  IVSVTX4 U2268 ( .A(n492), .Z(n3886) );
  B_ND2SVTX2 U2269 ( .A(n3667), .B(n3668), .Z(n3671) );
  IVSVTX4 U2270 ( .A(n993), .Z(n958) );
  IVSVTX4 U2271 ( .A(n2972), .Z(n1353) );
  AO7SVTX6 U2272 ( .A(n3452), .B(n3451), .C(n3450), .Z(n3521) );
  IVSVTX4 U2273 ( .A(n3089), .Z(n3090) );
  NR2SVTX4 U2274 ( .A(n2916), .B(n2915), .Z(n1502) );
  CTIVSVTX4 U2275 ( .A(n2881), .Z(n1041) );
  AO17ASVTX6 U2276 ( .A(n3282), .B(n1089), .C(n3067), .D(n2284), .Z(n2988) );
  CTIVSVTX2 U2277 ( .A(n2794), .Z(n2796) );
  IVSVTX2 U2278 ( .A(n1482), .Z(n1483) );
  IVSVTX2 U2279 ( .A(n1623), .Z(n871) );
  IVSVTX10 U2280 ( .A(n1484), .Z(n2789) );
  B_ND2SVTX2 U2281 ( .A(n621), .B(n3270), .Z(n2164) );
  IVSVTX4 U2282 ( .A(n3032), .Z(n1546) );
  CTIVSVTX2 U2283 ( .A(n2989), .Z(n2991) );
  IVSVTX8 U2284 ( .A(n619), .Z(n1089) );
  ND2ASVTX6 U2285 ( .A(n1642), .B(n2807), .Z(n914) );
  IVSVTX6 U2286 ( .A(n1759), .Z(n2944) );
  IVSVTX10 U2287 ( .A(n808), .Z(n1851) );
  IVSVTX8 U2288 ( .A(n814), .Z(n537) );
  ND2ASVTX6 U2289 ( .A(n1939), .B(n2149), .Z(n1826) );
  CTIVSVTX4 U2290 ( .A(n3460), .Z(n3083) );
  AO4ABSVTX6 U2291 ( .C(n2149), .D(n2148), .A(n3078), .B(n626), .Z(n2893) );
  IVSVTX2 U2292 ( .A(n1622), .Z(n1621) );
  IVSVTX6 U2293 ( .A(n1794), .Z(n613) );
  IVSVTX4 U2294 ( .A(n2918), .Z(n2903) );
  IVSVTX4 U2295 ( .A(n2138), .Z(n1912) );
  ND2SVTX2 U2296 ( .A(n2240), .B(n728), .Z(n1848) );
  IVSVTX6 U2297 ( .A(n2255), .Z(n2128) );
  CTBUFSVTX12 U2298 ( .A(n2370), .Z(n3270) );
  IVSVTX8 U2299 ( .A(n1647), .Z(n619) );
  AO7SVTX4 U2300 ( .A(n2993), .B(n3283), .C(n2353), .Z(n849) );
  IVSVTX10 U2301 ( .A(n2947), .Z(n3126) );
  IVSVTX10 U2302 ( .A(n3280), .Z(n2905) );
  ND2ASVTX4 U2303 ( .A(n1083), .B(n2704), .Z(n2318) );
  IVSVTX6 U2304 ( .A(n2784), .Z(n540) );
  IVSVTX8 U2305 ( .A(n1644), .Z(n1397) );
  IVSVTX10 U2306 ( .A(n1732), .Z(n1346) );
  BFSVTX12 U2307 ( .A(n1419), .Z(n541) );
  IVSVTX12 U2308 ( .A(n629), .Z(n545) );
  ND4ABSVTX6 U2309 ( .A(n1166), .B(n1677), .C(n2619), .D(n2330), .Z(n1252) );
  ND2SVTX4 U2310 ( .A(n682), .B(n2614), .Z(n681) );
  ND2SVTX4 U2311 ( .A(n1083), .B(n971), .Z(n1887) );
  AO20SVTX8 U2312 ( .A(n1605), .B(n902), .C(n2693), .D(n2694), .Z(n1604) );
  NR2SVTX6 U2313 ( .A(n1421), .B(n1774), .Z(n2331) );
  IVSVTX8 U2314 ( .A(n633), .Z(n548) );
  AO4SVTX4 U2315 ( .A(n2611), .B(n2612), .C(n1421), .D(n2613), .Z(n1420) );
  NR3SVTX4 U2316 ( .A(n2689), .B(n2690), .C(n634), .Z(n903) );
  ND2SVTX4 U2317 ( .A(n1576), .B(n2654), .Z(n1114) );
  IVSVTX2 U2318 ( .A(n2332), .Z(n2692) );
  IVSVTX10 U2319 ( .A(n2898), .Z(n549) );
  ND3SVTX6 U2320 ( .A(n1360), .B(n857), .C(n1022), .Z(n1230) );
  AO6CSVTX4 U2321 ( .A(n1772), .B(n1773), .C(n2312), .Z(n967) );
  IVSVTX4 U2322 ( .A(n1772), .Z(n2287) );
  ND2SVTX4 U2323 ( .A(n2503), .B(n1708), .Z(n2538) );
  ND2ASVTX4 U2324 ( .A(n635), .B(n513), .Z(n2659) );
  ND2ASVTX6 U2325 ( .A(n1564), .B(n2232), .Z(n2595) );
  IVSVTX10 U2326 ( .A(n1756), .Z(n1769) );
  NR3ABSVTX4 U2327 ( .A(n1568), .B(n861), .C(n2572), .Z(n1567) );
  IVSVTX8 U2328 ( .A(n2033), .Z(n2528) );
  ND2SVTX6 U2329 ( .A(n637), .B(n2133), .Z(n2177) );
  IVSVTX2 U2330 ( .A(n2588), .Z(n2589) );
  CTIVSVTX2 U2331 ( .A(n2698), .Z(n656) );
  NR2SVTX6 U2332 ( .A(num_i[30]), .B(num_i[31]), .Z(n2489) );
  NR2SVTX6 U2333 ( .A(num_i[11]), .B(num_i[10]), .Z(n2192) );
  CTIVSVTX4 U2334 ( .A(num_i[13]), .Z(n638) );
  IVSVTX4 U2335 ( .A(num_i[8]), .Z(n554) );
  AO6SVTX4 U2336 ( .A(n4306), .B(n1625), .C(n1731), .Z(n1624) );
  AO20SVTX4 U2337 ( .A(n1737), .B(n1736), .C(n1735), .D(n4271), .Z(n4275) );
  ENSVTX4 U2338 ( .A(n4307), .B(n4306), .Z(rslt_o[15]) );
  IVSVTX4 U2339 ( .A(n4274), .Z(n1735) );
  AO7SVTX4 U2340 ( .A(n4166), .B(n4207), .C(n1659), .Z(n1803) );
  ENSVTX4 U2341 ( .A(n2447), .B(n4218), .Z(rslt_o[10]) );
  IVSVTX2 U2342 ( .A(n4191), .Z(n1625) );
  AO6SVTX2 U2343 ( .A(n4301), .B(n4295), .C(n4297), .Z(n4227) );
  ENSVTX4 U2344 ( .A(n4233), .B(n4232), .Z(rslt_o[7]) );
  AO6SVTX2 U2345 ( .A(n4301), .B(n4242), .C(n4217), .Z(n4218) );
  ENSVTX4 U2346 ( .A(n4240), .B(n4239), .Z(rslt_o[8]) );
  F_AN2SVTX2 U2347 ( .A(n4148), .B(n4269), .Z(n4276) );
  AO7SVTX2 U2348 ( .A(n414), .B(n4245), .C(n4235), .Z(n4232) );
  AO7SVTX2 U2349 ( .A(n4238), .B(n4245), .C(n4237), .Z(n4239) );
  IVSVTX6 U2350 ( .A(n4196), .Z(n556) );
  AO7SVTX6 U2351 ( .A(n1014), .B(n4049), .C(n4048), .Z(n4220) );
  B_ND2SVTX2 U2352 ( .A(n4289), .B(n4288), .Z(n4292) );
  IVSVTX4 U2353 ( .A(n1464), .Z(n4277) );
  NR2SVTX6 U2354 ( .A(n939), .B(n935), .Z(n1716) );
  CTIVSVTX2 U2355 ( .A(n1720), .Z(n4226) );
  IVSVTX4 U2356 ( .A(n4278), .Z(n1008) );
  IVSVTX4 U2357 ( .A(n4086), .Z(n1467) );
  ND3SVTX4 U2358 ( .A(n1783), .B(n1782), .C(n4129), .Z(n1781) );
  B_ND2SVTX2 U2359 ( .A(n4254), .B(n4249), .Z(n4255) );
  B_ND2SVTX2 U2360 ( .A(n4263), .B(n797), .Z(n4264) );
  IVSVTX4 U2361 ( .A(n1402), .Z(n936) );
  ND2SVTX4 U2362 ( .A(n2235), .B(n1707), .Z(n1501) );
  NR4ABSVTX6 U2363 ( .A(n3197), .B(n3196), .C(n3195), .D(n3194), .Z(n3198) );
  IVSVTX2 U2364 ( .A(n2432), .Z(n2769) );
  ND2SVTX4 U2365 ( .A(n1414), .B(n1413), .Z(n934) );
  NR2SVTX6 U2366 ( .A(n2188), .B(n2186), .Z(n1845) );
  ND2SVTX4 U2367 ( .A(n4127), .B(n1778), .Z(n1782) );
  NR2SVTX2 U2368 ( .A(n4236), .B(n2383), .Z(n4237) );
  IVSVTX4 U2369 ( .A(n1411), .Z(n933) );
  ND3ASVTX6 U2370 ( .A(n1443), .B(n4164), .C(n1442), .Z(n1441) );
  B_ND2SVTX2 U2371 ( .A(n4168), .B(n2414), .Z(n4169) );
  IVSVTX2 U2372 ( .A(n4064), .Z(n1703) );
  ND4SVTX6 U2373 ( .A(n1628), .B(n940), .C(n1987), .D(n1392), .Z(n939) );
  AO3SVTX6 U2374 ( .A(n1896), .B(n4077), .C(n4076), .D(n4078), .Z(n4084) );
  AO6CSVTX6 U2375 ( .A(n1469), .B(n1468), .C(n2400), .Z(n916) );
  ND3SVTX4 U2376 ( .A(n751), .B(n986), .C(n750), .Z(n985) );
  ND2SVTX4 U2377 ( .A(n4131), .B(n4137), .Z(n1780) );
  ND2SVTX4 U2378 ( .A(n860), .B(n1073), .Z(n1072) );
  ND4ASVTX4 U2379 ( .A(n3249), .B(n3256), .C(n2041), .D(n3255), .Z(n2040) );
  ND2ASVTX4 U2380 ( .A(n4123), .B(n4178), .Z(n4127) );
  ND3SVTX4 U2381 ( .A(n1646), .B(n889), .C(n888), .Z(n1453) );
  ND3SVTX4 U2382 ( .A(n870), .B(n2021), .C(n2022), .Z(n2274) );
  ND3SVTX4 U2383 ( .A(n4091), .B(n529), .C(n3340), .Z(n1412) );
  IVSVTX2 U2384 ( .A(n1897), .Z(n747) );
  F_AN2SVTX2 U2385 ( .A(n2346), .B(n4091), .Z(n2414) );
  NR3ABSVTX6 U2386 ( .A(n3972), .B(n3701), .C(n1639), .Z(n2411) );
  AO8DSVTX4 U2387 ( .A(n3330), .B(n789), .C(n788), .D(n790), .Z(n1263) );
  AO7SVTX2 U2388 ( .A(n4161), .B(n4156), .C(n1911), .Z(n1443) );
  NR2SVTX4 U2389 ( .A(n3153), .B(n3152), .Z(n1645) );
  NR3SVTX4 U2390 ( .A(n3943), .B(n3942), .C(n905), .Z(n1184) );
  AO1SVTX4 U2391 ( .A(n483), .B(n3375), .C(n1862), .D(n2267), .Z(n987) );
  IVSVTX4 U2392 ( .A(n2085), .Z(n1278) );
  NR2ASVTX6 U2393 ( .A(n3221), .B(n2046), .Z(n2043) );
  ND2ASVTX4 U2394 ( .A(n1790), .B(n3144), .Z(n1667) );
  IVSVTX2 U2395 ( .A(n2386), .Z(n1476) );
  AO6SVTX4 U2396 ( .A(n3295), .B(n3296), .C(n1291), .Z(n940) );
  ND2SVTX4 U2397 ( .A(n4036), .B(n2311), .Z(n2310) );
  ND3ABSVTX6 U2398 ( .A(n493), .B(n2230), .C(n2444), .Z(n1081) );
  ND2SVTX4 U2399 ( .A(n2247), .B(n818), .Z(n723) );
  IVSVTX2 U2400 ( .A(n1172), .Z(n4061) );
  AO3CDSVTX4 U2401 ( .A(n2461), .B(n3228), .C(n3227), .D(n3226), .Z(n3233) );
  NR2SVTX4 U2402 ( .A(n1901), .B(n1849), .Z(n1897) );
  ND2SVTX4 U2403 ( .A(n615), .B(n4125), .Z(n1779) );
  ND3SVTX4 U2404 ( .A(n3329), .B(n3331), .C(n788), .Z(n1415) );
  CTIVSVTX2 U2405 ( .A(n4142), .Z(n4143) );
  AO7SVTX2 U2406 ( .A(n4040), .B(n4038), .C(n4037), .Z(n4045) );
  IVSVTX2 U2407 ( .A(n1429), .Z(n3158) );
  IVSVTX2 U2408 ( .A(n3218), .Z(n2173) );
  AO7SVTX4 U2409 ( .A(n3615), .B(n3614), .C(n3613), .Z(n3616) );
  AO7SVTX4 U2410 ( .A(n523), .B(n3297), .C(n2433), .Z(n1291) );
  IVSVTX2 U2411 ( .A(n3250), .Z(n2041) );
  ND4ABSVTX6 U2412 ( .A(n3582), .B(n3581), .C(n3580), .D(n3579), .Z(n3617) );
  ND2SVTX6 U2413 ( .A(n2135), .B(n3164), .Z(n2134) );
  IVSVTX2 U2414 ( .A(n3131), .Z(n2082) );
  NR3SVTX4 U2415 ( .A(n3339), .B(n3338), .C(n2113), .Z(n3340) );
  F_AN2SVTX2 U2416 ( .A(n4174), .B(n1715), .Z(n2440) );
  IVSVTX2 U2417 ( .A(n2278), .Z(n2021) );
  ND2SVTX4 U2418 ( .A(n3419), .B(n1900), .Z(n1849) );
  NR2SVTX4 U2419 ( .A(n1406), .B(n3319), .Z(n1405) );
  ND2SVTX4 U2420 ( .A(n2346), .B(n1715), .Z(n1157) );
  NR3SVTX4 U2421 ( .A(n4074), .B(n4073), .C(n4082), .Z(n4076) );
  ND4ABSVTX6 U2422 ( .A(n2291), .B(n3431), .C(n1100), .D(n1619), .Z(n818) );
  NR3SVTX6 U2423 ( .A(n2422), .B(n3968), .C(n1195), .Z(n1194) );
  ND2ASVTX4 U2424 ( .A(n3268), .B(n2096), .Z(n2095) );
  AO7SVTX4 U2425 ( .A(n3336), .B(n3335), .C(n865), .Z(n2278) );
  ND3SVTX4 U2426 ( .A(n1328), .B(n3337), .C(n514), .Z(n3338) );
  IVSVTX2 U2427 ( .A(n3567), .Z(n3582) );
  IVSVTX4 U2428 ( .A(n1880), .Z(n1879) );
  B_ND2SVTX2 U2429 ( .A(n3854), .B(n3188), .Z(n3189) );
  NR2SVTX2 U2430 ( .A(n3315), .B(n883), .Z(n3317) );
  ND2SVTX2 U2431 ( .A(n3575), .B(n1489), .Z(n3580) );
  AO20SVTX2 U2432 ( .A(n1983), .B(n4172), .C(n367), .D(n1422), .Z(n4183) );
  NR2SVTX4 U2433 ( .A(n1423), .B(n1424), .Z(n3825) );
  IVSVTX2 U2434 ( .A(n4065), .Z(n2218) );
  ND3SVTX4 U2435 ( .A(n2443), .B(n2396), .C(n3967), .Z(n1187) );
  IVSVTX2 U2436 ( .A(n3339), .Z(n3220) );
  ND3SVTX4 U2437 ( .A(n2350), .B(n1399), .C(n1398), .Z(n2174) );
  AO7NSVTX4 U2438 ( .A(n3877), .B(n1864), .C(n3876), .Z(n2444) );
  NR2ASVTX4 U2439 ( .A(n514), .B(n2425), .Z(n3221) );
  AN2SVTX2 U2440 ( .A(n3381), .B(n3854), .Z(n2271) );
  ND2SVTX6 U2441 ( .A(n1556), .B(n1555), .Z(n1557) );
  IVSVTX8 U2442 ( .A(n1550), .Z(n1715) );
  NR2ASVTX4 U2443 ( .A(n3613), .B(n3683), .Z(n1381) );
  NR2SVTX2 U2444 ( .A(n3181), .B(n3183), .Z(n2201) );
  IVSVTX2 U2445 ( .A(n887), .Z(n2160) );
  AO2SVTX4 U2446 ( .A(n445), .B(n4072), .C(n862), .D(n4071), .Z(n4082) );
  NR2SVTX2 U2447 ( .A(n3305), .B(n3302), .Z(n3304) );
  NR3SVTX6 U2448 ( .A(n1863), .B(n1260), .C(n3824), .Z(n1423) );
  ND2SVTX6 U2449 ( .A(n3235), .B(n3237), .Z(n1367) );
  NR2ASVTX4 U2450 ( .A(n3239), .B(n3230), .Z(n3227) );
  IVSVTX2 U2451 ( .A(n3750), .Z(n3752) );
  IVSVTX4 U2452 ( .A(n2233), .Z(n561) );
  IVSVTX2 U2453 ( .A(n3708), .Z(n3715) );
  IVSVTX2 U2454 ( .A(n3934), .Z(n1632) );
  ND2SVTX4 U2455 ( .A(n3961), .B(n3962), .Z(n3968) );
  AO6SVTX2 U2456 ( .A(n3361), .B(n3387), .C(n2273), .Z(n2272) );
  AO7SVTX6 U2457 ( .A(n3401), .B(n3397), .C(n2408), .Z(n1847) );
  NR3SVTX2 U2458 ( .A(n4093), .B(n3213), .C(n3211), .Z(n2410) );
  ND3SVTX4 U2459 ( .A(n927), .B(n3833), .C(n925), .Z(n754) );
  IVSVTX2 U2460 ( .A(n3387), .Z(n3363) );
  IVSVTX4 U2461 ( .A(n2451), .Z(n898) );
  IVSVTX2 U2462 ( .A(n3379), .Z(n1240) );
  AO7SVTX4 U2463 ( .A(n3206), .B(n3264), .C(n3205), .Z(n3208) );
  IVSVTX2 U2464 ( .A(n3380), .Z(n1602) );
  IVSVTX4 U2465 ( .A(n1135), .Z(n1134) );
  OR3SVTX4 U2466 ( .A(n3938), .B(n3937), .C(n3940), .Z(n3936) );
  NR2SVTX2 U2467 ( .A(n4073), .B(n3019), .Z(n1559) );
  IVSVTX4 U2468 ( .A(n1854), .Z(n1398) );
  NR2SVTX2 U2469 ( .A(n3578), .B(n3577), .Z(n711) );
  IVSVTX4 U2470 ( .A(n3789), .Z(n2202) );
  AO7SVTX4 U2471 ( .A(n3879), .B(n3877), .C(n3613), .Z(n2230) );
  IVSVTX4 U2472 ( .A(n1427), .Z(n1217) );
  NR2SVTX2 U2473 ( .A(n1289), .B(n4060), .Z(n4062) );
  ND2ASVTX4 U2474 ( .A(n3367), .B(n3307), .Z(n3306) );
  CTBUFSVTX12 U2475 ( .A(n2424), .Z(n4171) );
  CTIVSVTX2 U2476 ( .A(n3188), .Z(n3167) );
  AO7ASVTX6 U2477 ( .A(n3324), .B(n3264), .C(n3372), .Z(n2097) );
  NR2ASVTX4 U2478 ( .A(n3324), .B(n1635), .Z(n2099) );
  IVSVTX4 U2479 ( .A(n3234), .Z(n564) );
  ND2SVTX2 U2480 ( .A(n530), .B(n3360), .Z(n2273) );
  ND3SVTX4 U2481 ( .A(n3312), .B(n3246), .C(n3334), .Z(n3248) );
  IVSVTX2 U2482 ( .A(n2222), .Z(n1734) );
  IVSVTX4 U2483 ( .A(n3319), .Z(n565) );
  IVSVTX2 U2484 ( .A(n1725), .Z(n787) );
  ND2SVTX6 U2485 ( .A(n3965), .B(n744), .Z(n3266) );
  ND3SVTX4 U2486 ( .A(n831), .B(n2431), .C(n869), .Z(n3689) );
  F_ENSVTX2 U2487 ( .A(n3786), .B(n3785), .Z(n2109) );
  AO6ABSVTX4 U2488 ( .A(n3945), .B(n4006), .C(n697), .Z(n1340) );
  B_ND2SVTX2 U2489 ( .A(n4056), .B(n3229), .Z(n3232) );
  IVSVTX6 U2490 ( .A(n3792), .Z(n3929) );
  CTIVSVTX2 U2491 ( .A(n2425), .Z(n3258) );
  B_ND2SVTX2 U2492 ( .A(n4101), .B(n4100), .Z(n4103) );
  ND3SVTX4 U2493 ( .A(n3774), .B(n3773), .C(n1658), .Z(n3775) );
  CTIVSVTX4 U2494 ( .A(n2065), .Z(n2064) );
  IVSVTX2 U2495 ( .A(n3254), .Z(n1614) );
  NR2SVTX4 U2496 ( .A(n3427), .B(n3425), .Z(n3424) );
  IVSVTX6 U2497 ( .A(n2007), .Z(n3618) );
  IVSVTX2 U2498 ( .A(n3148), .Z(n2948) );
  IVSVTX4 U2499 ( .A(n2078), .Z(n1205) );
  ND2SVTX6 U2500 ( .A(n2325), .B(n2324), .Z(n3490) );
  AO7SVTX6 U2501 ( .A(n3332), .B(n3173), .C(n3245), .Z(n3184) );
  NR2SVTX4 U2502 ( .A(n3694), .B(n3695), .Z(n3696) );
  IVSVTX2 U2503 ( .A(n926), .Z(n3830) );
  IVSVTX4 U2504 ( .A(n1065), .Z(n1064) );
  IVSVTX2 U2505 ( .A(n534), .Z(n740) );
  ND3ASVTX6 U2506 ( .A(n3474), .B(n3558), .C(n3476), .Z(n1216) );
  CTIVSVTX4 U2507 ( .A(n2939), .Z(n1496) );
  IVSVTX2 U2508 ( .A(n3321), .Z(n3217) );
  ND2SVTX6 U2509 ( .A(n3690), .B(n1905), .Z(n1264) );
  IVSVTX4 U2510 ( .A(n2190), .Z(n2019) );
  NR2SVTX6 U2511 ( .A(n3585), .B(n3586), .Z(n2423) );
  ND2SVTX6 U2512 ( .A(n2066), .B(n1435), .Z(n710) );
  ND2SVTX6 U2513 ( .A(n2178), .B(n2824), .Z(n3924) );
  CTBUFSVTX4 U2514 ( .A(n4133), .Z(n775) );
  IVSVTX10 U2515 ( .A(n694), .Z(n2292) );
  AO7SVTX4 U2516 ( .A(n3870), .B(n1299), .C(n3871), .Z(n1425) );
  CTIVSVTX4 U2517 ( .A(n1511), .Z(n1512) );
  AO17ASVTX6 U2518 ( .A(n510), .B(n1146), .C(n505), .D(n1144), .Z(n1510) );
  IVSVTX2 U2519 ( .A(n1865), .Z(n1260) );
  OR2SVTX4 U2520 ( .A(n3374), .B(n3373), .Z(n3377) );
  B_ND2SVTX2 U2521 ( .A(n3707), .B(n3664), .Z(n3665) );
  IVSVTX4 U2522 ( .A(n3418), .Z(n881) );
  NR2ASVTX4 U2523 ( .A(n2190), .B(n1934), .Z(n1192) );
  CTBUFSVTX4 U2524 ( .A(n2336), .Z(n869) );
  IVSVTX2 U2525 ( .A(n3398), .Z(n1909) );
  IVSVTX6 U2526 ( .A(n3473), .Z(n3558) );
  ND2SVTX6 U2527 ( .A(n2153), .B(n2336), .Z(n3855) );
  IVSVTX4 U2528 ( .A(n3939), .Z(n4011) );
  IVSVTX2 U2529 ( .A(n3633), .Z(n3634) );
  AO6SVTX2 U2530 ( .A(n3624), .B(n2427), .C(n3598), .Z(n3599) );
  IVSVTX2 U2531 ( .A(n3823), .Z(n1865) );
  B_ND2SVTX2 U2532 ( .A(n3681), .B(n3808), .Z(n3682) );
  IVSVTX4 U2533 ( .A(n3511), .Z(n3512) );
  B_ND2SVTX2 U2534 ( .A(n3545), .B(n2450), .Z(n3546) );
  NR2ASVTX4 U2535 ( .A(n3704), .B(n3707), .Z(n3711) );
  IVSVTX4 U2536 ( .A(n1934), .Z(n1935) );
  ND2ASVTX4 U2537 ( .A(n1004), .B(n2809), .Z(n3999) );
  AO7ABSVTX4 U2538 ( .A(n3841), .B(n1305), .C(n1663), .Z(n2338) );
  IVSVTX6 U2539 ( .A(n3219), .Z(n573) );
  ND2SVTX6 U2540 ( .A(n2715), .B(n2716), .Z(n2260) );
  IVSVTX6 U2541 ( .A(n1516), .Z(n1884) );
  ND2SVTX6 U2542 ( .A(n2163), .B(n2162), .Z(n2939) );
  ND2SVTX4 U2543 ( .A(n3291), .B(n3888), .Z(n1500) );
  B_ND2SVTX2 U2544 ( .A(n3612), .B(n3681), .Z(n3609) );
  ND2SVTX6 U2545 ( .A(n3093), .B(n1238), .Z(n3087) );
  CTIVSVTX4 U2546 ( .A(n4001), .Z(n575) );
  AO7SVTX6 U2547 ( .A(n1516), .B(n3853), .C(n3763), .Z(n3418) );
  AO3SVTX6 U2548 ( .A(n3422), .B(n1079), .C(n3973), .D(n3420), .Z(n3203) );
  ND2SVTX4 U2549 ( .A(n3956), .B(n3955), .Z(n3969) );
  B_ND2SVTX2 U2550 ( .A(n2950), .B(n2951), .Z(n3151) );
  CTIVSVTX2 U2551 ( .A(n3949), .Z(n3954) );
  CTAN2BSVTX4 U2552 ( .A(n3458), .B(n3461), .Z(n3472) );
  IVSVTX2 U2553 ( .A(n923), .Z(n922) );
  ND2SVTX4 U2554 ( .A(n2895), .B(n3772), .Z(n2153) );
  NR2SVTX6 U2555 ( .A(n811), .B(n810), .Z(n2895) );
  ND2SVTX6 U2556 ( .A(n1237), .B(n1236), .Z(n1238) );
  AN2SVTX4 U2557 ( .A(n3684), .B(n3597), .Z(n2427) );
  CTIVSVTX2 U2558 ( .A(n4145), .Z(n578) );
  CTIVSVTX4 U2559 ( .A(n3224), .Z(n580) );
  IVSVTX2 U2560 ( .A(n3461), .Z(n803) );
  ND3SVTX4 U2561 ( .A(n3980), .B(n3411), .C(n3764), .Z(n2000) );
  IVSVTX2 U2562 ( .A(n3393), .Z(n859) );
  AO7SVTX4 U2563 ( .A(n1177), .B(n2912), .C(n3412), .Z(n1220) );
  AO17ASVTX6 U2564 ( .A(n1251), .B(n2945), .C(n2807), .D(n1256), .Z(n2866) );
  ND2SVTX6 U2565 ( .A(n3702), .B(n2371), .Z(n3712) );
  AO1CDSVTX6 U2566 ( .A(n1962), .B(n3675), .C(n1960), .D(n3667), .Z(n3640) );
  IVSVTX4 U2567 ( .A(n3584), .Z(n3587) );
  NR2SVTX6 U2568 ( .A(n2963), .B(n2962), .Z(n3374) );
  AO7SVTX6 U2569 ( .A(n3603), .B(n3290), .C(n3636), .Z(n3888) );
  ND2SVTX6 U2570 ( .A(n2963), .B(n2962), .Z(n3372) );
  B_ND2SVTX2 U2571 ( .A(n3367), .B(n3366), .Z(n3381) );
  CTIVSVTX2 U2572 ( .A(n3137), .Z(n3139) );
  AO17ASVTX6 U2573 ( .A(n3435), .B(n1959), .C(n3434), .D(n1958), .Z(n3641) );
  CTBUFSVTX4 U2574 ( .A(n3393), .Z(n4030) );
  AO7ABSVTX4 U2575 ( .A(n2344), .B(n1088), .C(n896), .Z(n695) );
  IVSVTX4 U2576 ( .A(n3093), .Z(n3812) );
  CTIVSVTX2 U2577 ( .A(n3036), .Z(n3033) );
  B_ND2SVTX2 U2578 ( .A(n3125), .B(n3111), .Z(n3030) );
  IVSVTX2 U2579 ( .A(n2328), .Z(n2327) );
  CTIVSVTX4 U2580 ( .A(n4140), .Z(n589) );
  NR2ASVTX4 U2581 ( .A(n3126), .B(n3125), .Z(n3026) );
  ND2SVTX6 U2582 ( .A(n1714), .B(n1985), .Z(n3933) );
  IVSVTX4 U2583 ( .A(n3638), .Z(n3290) );
  B_ND2SVTX2 U2584 ( .A(n2412), .B(n2928), .Z(n3137) );
  AO7ABSVTX4 U2585 ( .A(n1851), .B(n1526), .C(n2060), .Z(n2329) );
  ND2SVTX4 U2586 ( .A(n3691), .B(n1327), .Z(n1980) );
  IVSVTX4 U2587 ( .A(n3661), .Z(n1513) );
  IVSVTX4 U2588 ( .A(n3040), .Z(n773) );
  IVSVTX4 U2589 ( .A(n3095), .Z(n1237) );
  IVSVTX4 U2590 ( .A(n2951), .Z(n2952) );
  F_ND2ASVTX2 U2591 ( .A(n1825), .B(n3672), .Z(n3436) );
  NR2SVTX4 U2592 ( .A(n3009), .B(n3008), .Z(n1077) );
  F_ND2SVTX1 U2593 ( .A(n3386), .B(n3385), .Z(n3388) );
  AO7SVTX6 U2594 ( .A(n3704), .B(n2894), .C(n3702), .Z(n3416) );
  CTIVSVTX4 U2595 ( .A(n2795), .Z(n591) );
  IVSVTX4 U2596 ( .A(n510), .Z(n1063) );
  IVSVTX4 U2597 ( .A(n2781), .Z(n2779) );
  ND2SVTX6 U2598 ( .A(n2169), .B(n1437), .Z(n1450) );
  AO17CSVTX6 U2599 ( .A(n3519), .B(n3521), .C(n3508), .D(n794), .Z(n1506) );
  ND2SVTX6 U2600 ( .A(n2872), .B(n2873), .Z(n3367) );
  ND2SVTX6 U2601 ( .A(n1434), .B(n1433), .Z(n2862) );
  CTIVSVTX2 U2602 ( .A(n3626), .Z(n885) );
  NR2ASVTX4 U2603 ( .A(n2358), .B(n3414), .Z(n3765) );
  ND2ASVTX6 U2604 ( .A(n757), .B(n1344), .Z(n3813) );
  CTIVSVTX2 U2605 ( .A(n2930), .Z(n2931) );
  B_ND2SVTX2 U2606 ( .A(n4006), .B(n3945), .Z(n3938) );
  CTIVSVTX4 U2607 ( .A(n2894), .Z(n2371) );
  IVSVTX2 U2608 ( .A(n3858), .Z(n592) );
  IVSVTX2 U2609 ( .A(n3454), .Z(n2459) );
  NR2SVTX6 U2610 ( .A(n3504), .B(n3503), .Z(n3080) );
  ND2ASVTX6 U2611 ( .A(n2798), .B(n2800), .Z(n2933) );
  B_ND2SVTX2 U2612 ( .A(n615), .B(n1790), .Z(n3036) );
  ND2SVTX6 U2613 ( .A(n2821), .B(n2823), .Z(n2120) );
  IVSVTX2 U2614 ( .A(n1368), .Z(n757) );
  IVSVTX4 U2615 ( .A(n2823), .Z(n1019) );
  IVSVTX6 U2616 ( .A(n1521), .Z(n1369) );
  IVSVTX2 U2617 ( .A(n3025), .Z(n3029) );
  ND2SVTX4 U2618 ( .A(n2847), .B(n2191), .Z(n1433) );
  ND2SVTX6 U2619 ( .A(n1979), .B(n1771), .Z(n1327) );
  NR2SVTX6 U2620 ( .A(n3554), .B(n1261), .Z(n794) );
  CTBUFSVTX4 U2621 ( .A(n3625), .Z(n1665) );
  CTIVSVTX2 U2622 ( .A(n930), .Z(n596) );
  ND2SVTX4 U2623 ( .A(n408), .B(n3570), .Z(n2152) );
  AO7SVTX2 U2624 ( .A(n4006), .B(n4007), .C(n2301), .Z(n4008) );
  IVSVTX2 U2625 ( .A(n2388), .Z(n1984) );
  ND2SVTX6 U2626 ( .A(n2889), .B(n2890), .Z(n3552) );
  AO6SVTX2 U2627 ( .A(n3935), .B(n2157), .C(n4005), .Z(n2156) );
  B_ND2SVTX2 U2628 ( .A(n3887), .B(n3886), .Z(n3891) );
  ND2SVTX4 U2629 ( .A(n2814), .B(n2813), .Z(n2170) );
  ND2SVTX4 U2630 ( .A(n2960), .B(n2961), .Z(n3267) );
  B_ND2SVTX2 U2631 ( .A(n3122), .B(n1254), .Z(n2958) );
  IVSVTX4 U2632 ( .A(n1809), .Z(n1808) );
  ND2ASVTX6 U2633 ( .A(n3286), .B(n3285), .Z(n3433) );
  IVSVTX6 U2634 ( .A(n2297), .Z(n598) );
  IVSVTX4 U2635 ( .A(n3011), .Z(n1080) );
  IVSVTX4 U2636 ( .A(n2911), .Z(n1204) );
  IVSVTX4 U2637 ( .A(n3959), .Z(n601) );
  IVSVTX4 U2638 ( .A(n3827), .Z(n602) );
  IVSVTX4 U2639 ( .A(n3046), .Z(n3042) );
  IVSVTX2 U2640 ( .A(n3459), .Z(n802) );
  IVSVTX6 U2641 ( .A(n3957), .Z(n1655) );
  IVSVTX2 U2642 ( .A(n3077), .Z(n3086) );
  F_IVSVTX1 U2643 ( .A(n3749), .Z(n3783) );
  IVSVTX4 U2644 ( .A(n2999), .Z(n732) );
  F_ND2ASVTX2 U2645 ( .A(n942), .B(n2348), .Z(n3358) );
  ND2SVTX6 U2646 ( .A(n703), .B(n2972), .Z(n3691) );
  IVSVTX2 U2647 ( .A(n2051), .Z(n2049) );
  IVSVTX2 U2648 ( .A(n4004), .Z(n2157) );
  B_ND2SVTX2 U2649 ( .A(n3494), .B(n3493), .Z(n3497) );
  CTBUFSVTX12 U2650 ( .A(n2789), .Z(n3014) );
  IVSVTX2 U2651 ( .A(n2727), .Z(n1650) );
  B_ND2SVTX2 U2652 ( .A(n652), .B(n3122), .Z(n2871) );
  ND2SVTX4 U2653 ( .A(n1851), .B(n1151), .Z(n1815) );
  OR2SVTX6 U2654 ( .A(n814), .B(n1892), .Z(n3098) );
  AO7SVTX4 U2655 ( .A(n1223), .B(n1791), .C(n1743), .Z(n1595) );
  IVSVTX2 U2656 ( .A(n3668), .Z(n1964) );
  ND2ASVTX6 U2657 ( .A(n728), .B(n1208), .Z(n1207) );
  CTIVSVTX4 U2658 ( .A(n2998), .Z(n605) );
  IVSVTX10 U2659 ( .A(n541), .Z(n1791) );
  AO7SVTX4 U2660 ( .A(n1972), .B(n2141), .C(n704), .Z(n703) );
  IVSVTX4 U2661 ( .A(n2878), .Z(n607) );
  ND2ASVTX6 U2662 ( .A(n2989), .B(n2990), .Z(n3522) );
  ND2ASVTX4 U2663 ( .A(n2760), .B(n1149), .Z(n2749) );
  IVSVTX4 U2664 ( .A(n3126), .Z(n611) );
  B_ND2SVTX2 U2665 ( .A(n728), .B(n503), .Z(n2460) );
  IVSVTX4 U2666 ( .A(n3477), .Z(n614) );
  ND2SVTX6 U2667 ( .A(n1882), .B(n3282), .Z(n3668) );
  ND2ASVTX6 U2668 ( .A(n2576), .B(n2703), .Z(n1853) );
  F_EOSVTX2 U2669 ( .A(n1347), .B(n942), .Z(n941) );
  ND2SVTX6 U2670 ( .A(n2319), .B(n2318), .Z(n1484) );
  ND2SVTX6 U2671 ( .A(n2888), .B(n911), .Z(n677) );
  IVSVTX10 U2672 ( .A(n839), .Z(n3273) );
  IVSVTX12 U2673 ( .A(n2370), .Z(n617) );
  IVSVTX6 U2674 ( .A(n2947), .Z(n618) );
  ND2SVTX4 U2675 ( .A(n548), .B(n2707), .Z(n1579) );
  ND2SVTX4 U2676 ( .A(n548), .B(n2707), .Z(n1570) );
  ND2SVTX6 U2677 ( .A(n2641), .B(n2640), .Z(n1142) );
  IVSVTX12 U2678 ( .A(n1419), .Z(n620) );
  IVSVTX4 U2679 ( .A(n518), .Z(n621) );
  BFSVTX12 U2680 ( .A(n2784), .Z(n622) );
  ND2SVTX6 U2681 ( .A(n947), .B(n945), .Z(n839) );
  ND3SVTX4 U2682 ( .A(n2839), .B(n2305), .C(n2307), .Z(n2701) );
  IVSVTX12 U2683 ( .A(n2971), .Z(n625) );
  AN3CSVTX6 U2684 ( .A(n2621), .B(n2384), .C(n1701), .Z(n2752) );
  CTBUFSVTX8 U2685 ( .A(n1748), .Z(n626) );
  IVSVTX4 U2686 ( .A(n2143), .Z(n1859) );
  IVSVTX10 U2687 ( .A(n1265), .Z(n1268) );
  IVSVTX8 U2688 ( .A(n547), .Z(n627) );
  ND2SVTX6 U2689 ( .A(n1165), .B(n1044), .Z(n1265) );
  IVSVTX8 U2690 ( .A(n836), .Z(n628) );
  CTBUFSVTX4 U2691 ( .A(n1178), .Z(n1721) );
  IVSVTX4 U2692 ( .A(n1604), .Z(n2702) );
  IVSVTX2 U2693 ( .A(n1860), .Z(n2384) );
  ND2SVTX6 U2694 ( .A(n2568), .B(n1724), .Z(n2059) );
  ND2SVTX6 U2695 ( .A(n2183), .B(n951), .Z(n2550) );
  NR2SVTX4 U2696 ( .A(n1687), .B(n2331), .Z(n2330) );
  IVSVTX8 U2697 ( .A(n899), .Z(n629) );
  IVSVTX4 U2698 ( .A(n2760), .Z(n630) );
  ND2SVTX4 U2699 ( .A(n1772), .B(n1514), .Z(n2568) );
  NR2ASVTX6 U2700 ( .A(n2449), .B(n676), .Z(n2668) );
  IVSVTX12 U2701 ( .A(n1166), .Z(n631) );
  IVSVTX4 U2702 ( .A(n884), .Z(n834) );
  ND3SVTX4 U2703 ( .A(n2684), .B(n1656), .C(n2683), .Z(n2693) );
  ND2SVTX6 U2704 ( .A(n1656), .B(n2686), .Z(n1055) );
  IVSVTX4 U2705 ( .A(n2609), .Z(n1153) );
  IVSVTX2 U2706 ( .A(n2699), .Z(n1648) );
  NR2ASVTX4 U2707 ( .A(n920), .B(n2697), .Z(n2685) );
  NR2ASVTX6 U2708 ( .A(n1773), .B(n2287), .Z(n1971) );
  IVSVTX12 U2709 ( .A(n1107), .Z(n2636) );
  ND2SVTX4 U2710 ( .A(n2503), .B(n1037), .Z(n1038) );
  CTBUFSVTX12 U2711 ( .A(n2126), .Z(n895) );
  OR2SVTX2 U2712 ( .A(n2625), .B(n2364), .Z(n2449) );
  AO7SVTX6 U2713 ( .A(n912), .B(n963), .C(n2494), .Z(n1584) );
  IVSVTX4 U2714 ( .A(n2530), .Z(n2281) );
  AO7SVTX6 U2715 ( .A(n2519), .B(n2520), .C(n550), .Z(n2521) );
  ND3SVTX8 U2716 ( .A(n674), .B(n672), .C(n673), .Z(n2246) );
  ND2SVTX2 U2717 ( .A(n2488), .B(n963), .Z(n2127) );
  ND3SVTX4 U2718 ( .A(n2193), .B(n2145), .C(n2192), .Z(n2144) );
  ND2SVTX6 U2719 ( .A(n2498), .B(n2377), .Z(n1586) );
  F_ND2SVTX1 U2720 ( .A(num_i[3]), .B(n1744), .Z(n2625) );
  IVSVTX6 U2721 ( .A(n1410), .Z(n912) );
  ND3SVTX4 U2722 ( .A(num_i[7]), .B(n553), .C(n554), .Z(n2209) );
  CTBUFSVTX2 U2723 ( .A(num_i[10]), .Z(n2658) );
  CTBUFSVTX2 U2724 ( .A(num_i[11]), .Z(n2624) );
  NR2SVTX6 U2725 ( .A(num_i[5]), .B(num_i[7]), .Z(n1811) );
  NR2SVTX6 U2726 ( .A(num_i[4]), .B(num_i[6]), .Z(n1812) );
  IVSVTX4 U2727 ( .A(n451), .Z(n2671) );
  IVSVTX2 U2728 ( .A(num_i[2]), .Z(n2507) );
  CTBUFSVTX2 U2729 ( .A(num_i[6]), .Z(n920) );
  IVSVTX8 U2730 ( .A(num_i[27]), .Z(n639) );
  ND3ABSVTX8 U2731 ( .A(n3734), .B(n3733), .C(n3908), .Z(n641) );
  NR4ABCSVTX8 U2732 ( .A(n3972), .B(n3762), .C(n3761), .D(n641), .Z(n1890) );
  ND2SVTX4 U2733 ( .A(n566), .B(n641), .Z(n4293) );
  ND2ASVTX8 U2734 ( .A(n2222), .B(n3299), .Z(n642) );
  ND3SVTX6 U2735 ( .A(n642), .B(n558), .C(n1715), .Z(n767) );
  AO17SVTX4 U2736 ( .A(n642), .B(n559), .C(n467), .D(n2160), .Z(n1439) );
  AO4SVTX8 U2737 ( .A(n2806), .B(n2902), .C(n1287), .D(n706), .Z(n836) );
  AO7SVTX8 U2738 ( .A(n738), .B(n966), .C(n737), .Z(n706) );
  ND3SVTX8 U2739 ( .A(n2649), .B(n2650), .C(n2648), .Z(n2806) );
  NR2SVTX8 U2740 ( .A(n844), .B(n2172), .Z(n793) );
  ND3SVTX8 U2741 ( .A(n2050), .B(n2830), .C(n644), .Z(n844) );
  ND2SVTX8 U2742 ( .A(n2829), .B(n3839), .Z(n644) );
  IVSVTX4 U2743 ( .A(n645), .Z(n2672) );
  ND2SVTX6 U2744 ( .A(n1107), .B(n512), .Z(n2266) );
  IVSVTX4 U2745 ( .A(n647), .Z(n1875) );
  ND2ASVTX8 U2746 ( .A(n504), .B(n1533), .Z(n647) );
  ND3SVTX8 U2747 ( .A(n3021), .B(n660), .C(n2119), .Z(n1021) );
  IVSVTX4 U2748 ( .A(n2652), .Z(n2256) );
  ND2SVTX4 U2749 ( .A(n1233), .B(n2036), .Z(n707) );
  AO7SVTX6 U2750 ( .A(n2653), .B(n403), .C(n549), .Z(n649) );
  IVSVTX4 U2751 ( .A(n2258), .Z(n2653) );
  ND3ASVTX8 U2752 ( .A(n847), .B(n1015), .C(n1106), .Z(n1117) );
  IVSVTX12 U2753 ( .A(n651), .Z(n686) );
  ND2SVTX6 U2754 ( .A(n692), .B(n685), .Z(n651) );
  CTBUFSVTX2 U2755 ( .A(n3273), .Z(n652) );
  EN3SVTX8 U2756 ( .A(n2375), .B(n3273), .C(n2905), .Z(n2979) );
  IVSVTX4 U2757 ( .A(n2232), .Z(n2231) );
  NR2SVTX4 U2758 ( .A(n655), .B(n653), .Z(n886) );
  ND2ASVTX8 U2759 ( .A(n2491), .B(n654), .Z(n1219) );
  IVSVTX4 U2760 ( .A(n2551), .Z(n2491) );
  NR2SVTX4 U2761 ( .A(n658), .B(n666), .Z(n1913) );
  IVSVTX4 U2762 ( .A(n686), .Z(n691) );
  IVSVTX4 U2763 ( .A(n683), .Z(n659) );
  ND3SVTX8 U2764 ( .A(n1867), .B(n2726), .C(n1868), .Z(n660) );
  ND3ABSVTX8 U2765 ( .A(n1697), .B(n844), .C(n661), .Z(n3735) );
  AO20CSVTX8 U2766 ( .A(n3622), .B(n661), .C(n3623), .D(n4073), .Z(n3652) );
  ND3SVTX8 U2767 ( .A(n637), .B(n663), .C(n662), .Z(n2525) );
  NR2SVTX6 U2768 ( .A(num_i[28]), .B(num_i[24]), .Z(n662) );
  NR2SVTX6 U2769 ( .A(num_i[17]), .B(num_i[26]), .Z(n663) );
  AO7SVTX8 U2770 ( .A(n2314), .B(n665), .C(n2243), .Z(n2155) );
  IVSVTX4 U2771 ( .A(n669), .Z(n762) );
  NR2SVTX4 U2772 ( .A(n508), .B(n669), .Z(n668) );
  ND3ASVTX6 U2773 ( .A(n2387), .B(n2142), .C(n2288), .Z(n669) );
  ND2SVTX4 U2774 ( .A(n2718), .B(n1650), .Z(n3021) );
  F_EOSVTX2 U2775 ( .A(n3454), .B(n671), .Z(n670) );
  ND2SVTX4 U2776 ( .A(n1128), .B(n3524), .Z(n671) );
  ND4ASVTX6 U2777 ( .A(n2512), .B(n673), .C(n672), .D(n674), .Z(n690) );
  NR2ASVTX8 U2778 ( .A(n2497), .B(n2033), .Z(n674) );
  AO5ASVTX8 U2779 ( .B(n2240), .A(n1025), .C(n677), .Z(n716) );
  EN3SVTX8 U2780 ( .A(n2887), .B(n677), .C(n1089), .Z(n1087) );
  NR2SVTX4 U2781 ( .A(n3189), .B(n678), .Z(n3195) );
  ND2SVTX4 U2782 ( .A(n1270), .B(n3303), .Z(n678) );
  AN2SVTX8 U2783 ( .A(n2061), .B(n1246), .Z(n3303) );
  ND2SVTX8 U2784 ( .A(n3690), .B(n2336), .Z(n679) );
  ND2SVTX6 U2785 ( .A(n3983), .B(n679), .Z(n3732) );
  ND2SVTX4 U2786 ( .A(n679), .B(n1503), .Z(n1900) );
  ND2ASVTX8 U2787 ( .A(n1026), .B(n2322), .Z(n2641) );
  BFSVTX6 U2788 ( .A(n545), .Z(n687) );
  ND2ASVTX8 U2789 ( .A(n688), .B(n2882), .Z(n2884) );
  NR3SVTX8 U2790 ( .A(n1166), .B(n2059), .C(n693), .Z(n1418) );
  CTBUFSVTX12 U2791 ( .A(n3673), .Z(n697) );
  ND2SVTX4 U2792 ( .A(n3522), .B(n3588), .Z(n699) );
  NR2SVTX4 U2793 ( .A(n3673), .B(n702), .Z(n701) );
  ND2ASVTX8 U2794 ( .A(n703), .B(n1353), .Z(n3583) );
  ND2SVTX4 U2795 ( .A(n2971), .B(n1030), .Z(n704) );
  IVSVTX8 U2796 ( .A(n705), .Z(n3802) );
  ND2SVTX8 U2797 ( .A(n2360), .B(n3796), .Z(n705) );
  IVSVTX4 U2798 ( .A(n706), .Z(n971) );
  ND2SVTX4 U2799 ( .A(n680), .B(n706), .Z(n1528) );
  IVSVTX4 U2800 ( .A(n708), .Z(n3816) );
  NR2SVTX4 U2801 ( .A(n3607), .B(n3606), .Z(n708) );
  ND2ASVTX8 U2802 ( .A(n3606), .B(n3608), .Z(n3681) );
  ND2SVTX8 U2803 ( .A(n2125), .B(n2662), .Z(n798) );
  ND2SVTX8 U2804 ( .A(n1127), .B(n2279), .Z(n2662) );
  ND3SVTX8 U2805 ( .A(n713), .B(n3660), .C(n710), .Z(n1765) );
  ND2SVTX2 U2806 ( .A(n713), .B(n710), .Z(n796) );
  AO20SVTX8 U2807 ( .A(n1657), .B(n712), .C(n3659), .D(n2439), .Z(n1379) );
  IVSVTX4 U2808 ( .A(n1489), .Z(n712) );
  ND2ASVTX8 U2809 ( .A(n1450), .B(n1436), .Z(n713) );
  EO3SVTX8 U2810 ( .A(n538), .B(n716), .C(n2834), .Z(n1085) );
  EO3SVTX8 U2811 ( .A(n544), .B(n1685), .C(n1030), .Z(n2834) );
  AO7ABSVTX6 U2812 ( .A(n2887), .B(n684), .C(n2832), .Z(n2844) );
  ND2ASVTX8 U2813 ( .A(n3570), .B(n3443), .Z(n2006) );
  AO7ABSVTX4 U2814 ( .A(n3079), .B(n1149), .C(n714), .Z(n3570) );
  IVSVTX4 U2815 ( .A(n3065), .Z(n1149) );
  ND3SVTX8 U2816 ( .A(n3620), .B(n3618), .C(n3619), .Z(n715) );
  NR3ABSVTX8 U2817 ( .A(n2360), .B(n715), .C(n4023), .Z(n2197) );
  IVSVTX4 U2818 ( .A(n716), .Z(n1058) );
  ND3SVTX8 U2819 ( .A(n1532), .B(n1953), .C(n527), .Z(n3907) );
  AO7SVTX6 U2820 ( .A(n4250), .B(n720), .C(n1093), .Z(n724) );
  AO7SVTX6 U2821 ( .A(n719), .B(n718), .C(n717), .Z(n1093) );
  ND2SVTX4 U2822 ( .A(n856), .B(n722), .Z(n718) );
  NR2SVTX6 U2823 ( .A(n2250), .B(n1102), .Z(n721) );
  IVSVTX4 U2824 ( .A(n724), .Z(n3562) );
  CTBUFSVTX2 U2825 ( .A(n2540), .Z(n725) );
  NR2SVTX8 U2826 ( .A(n726), .B(n2177), .Z(n2540) );
  ND2SVTX8 U2827 ( .A(n639), .B(n640), .Z(n726) );
  IVSVTX4 U2828 ( .A(n726), .Z(n2481) );
  NR2ASVTX6 U2829 ( .A(n1551), .B(n804), .Z(n3071) );
  NR2SVTX8 U2830 ( .A(n545), .B(n798), .Z(n730) );
  ND2SVTX6 U2831 ( .A(n2636), .B(n2661), .Z(n1997) );
  ND2SVTX8 U2832 ( .A(n631), .B(n1178), .Z(n2321) );
  AO1CDSVTX8 U2833 ( .A(n1202), .B(n4271), .C(n3109), .D(n4148), .Z(n4207) );
  ND3SVTX6 U2834 ( .A(n3781), .B(n2073), .C(n3780), .Z(n731) );
  ND3SVTX8 U2835 ( .A(n1081), .B(n867), .C(n809), .Z(n829) );
  ND2ASVTX8 U2836 ( .A(n605), .B(n732), .Z(n3428) );
  NR2SVTX4 U2837 ( .A(n585), .B(n907), .Z(n3731) );
  ND2SVTX4 U2838 ( .A(n1045), .B(n1124), .Z(n1044) );
  AO7ABSVTX4 U2839 ( .A(n1972), .B(n2129), .C(n1836), .Z(n1368) );
  EO3SVTX8 U2840 ( .A(n686), .B(n2176), .C(n3068), .Z(n2995) );
  ND2SVTX4 U2841 ( .A(n2334), .B(n2902), .Z(n1052) );
  IVSVTX4 U2842 ( .A(n4219), .Z(n4029) );
  AO17CSVTX8 U2843 ( .A(n1023), .B(n2651), .C(n965), .D(n1060), .Z(n737) );
  EO3SVTX8 U2844 ( .A(n1481), .B(n997), .C(n959), .Z(n3621) );
  ND3ABSVTX6 U2845 ( .A(n1329), .B(n844), .C(n2171), .Z(n1597) );
  ND2SVTX4 U2846 ( .A(n476), .B(n4138), .Z(n1109) );
  NR2SVTX6 U2847 ( .A(n2496), .B(n2495), .Z(n1583) );
  F_ND3SVTX2 U2848 ( .A(n4032), .B(n3187), .C(n3186), .Z(n3196) );
  AO7SVTX6 U2849 ( .A(n4208), .B(n4207), .C(n1599), .Z(n4209) );
  BFSVTX1 U2850 ( .A(n1295), .Z(n741) );
  AO2SVTX4 U2851 ( .A(n2610), .B(n1576), .C(n1580), .D(n549), .Z(n2057) );
  ND2SVTX4 U2852 ( .A(n533), .B(n743), .Z(n2311) );
  ND2SVTX4 U2853 ( .A(n1718), .B(n3789), .Z(n743) );
  NR2ASVTX6 U2854 ( .A(n1766), .B(n1633), .Z(n3530) );
  AO7SVTX8 U2855 ( .A(n1003), .B(n970), .C(n2679), .Z(n2353) );
  ND3SVTX8 U2856 ( .A(n1350), .B(n2175), .C(n2038), .Z(n1349) );
  IVSVTX4 U2857 ( .A(n1352), .Z(n746) );
  NR2SVTX8 U2858 ( .A(n1914), .B(n4215), .Z(n4295) );
  ND3SVTX6 U2859 ( .A(n1968), .B(n909), .C(n908), .Z(n809) );
  ND2SVTX4 U2860 ( .A(n2326), .B(n1901), .Z(n749) );
  ND4SVTX6 U2861 ( .A(n1715), .B(n2346), .C(n4091), .D(n559), .Z(n4137) );
  IVSVTX10 U2862 ( .A(n686), .Z(n3067) );
  AO7ABSVTX8 U2863 ( .A(n3558), .B(n3466), .C(n648), .Z(n3467) );
  IVSVTX12 U2864 ( .A(n2570), .Z(n2561) );
  IVSVTX12 U2865 ( .A(n1142), .Z(n808) );
  NR2SVTX8 U2866 ( .A(n1076), .B(n1069), .Z(n4147) );
  IVSVTX4 U2867 ( .A(n1285), .Z(n1284) );
  ND2SVTX4 U2868 ( .A(n2370), .B(n1851), .Z(n3099) );
  IVSVTX8 U2869 ( .A(n562), .Z(n1235) );
  NR3ABSVTX8 U2870 ( .A(n3788), .B(n3740), .C(n4032), .Z(n3758) );
  EN3SVTX8 U2871 ( .A(n1647), .B(n1644), .C(n1764), .Z(n3088) );
  ND2SVTX4 U2872 ( .A(n1240), .B(n1241), .Z(n750) );
  ND2SVTX4 U2873 ( .A(n2271), .B(n4058), .Z(n751) );
  IVSVTX4 U2874 ( .A(n2066), .Z(n752) );
  AO5SVTX6 U2875 ( .A(n1526), .B(n1089), .C(n1889), .Z(n2973) );
  AO7SVTX6 U2876 ( .A(n3871), .B(n3812), .C(n3813), .Z(n2203) );
  IVSVTX8 U2877 ( .A(n847), .Z(n2620) );
  ND3ABSVTX8 U2878 ( .A(n635), .B(n2582), .C(n1544), .Z(n2501) );
  AO7SVTX8 U2879 ( .A(n3568), .B(n758), .C(n3565), .Z(n3162) );
  ND2SVTX4 U2880 ( .A(n2863), .B(n2864), .Z(n3565) );
  ND2ASVTX8 U2881 ( .A(n2015), .B(n2016), .Z(n3564) );
  ND2ASVTX8 U2882 ( .A(n2852), .B(n2851), .Z(n3566) );
  EO3SVTX8 U2883 ( .A(n1973), .B(n2854), .C(n2138), .Z(n2372) );
  IVSVTX4 U2884 ( .A(n2237), .Z(n2863) );
  EO3SVTX8 U2885 ( .A(n2858), .B(n1975), .C(n800), .Z(n2864) );
  IVSVTX4 U2886 ( .A(n914), .Z(n759) );
  ND3SVTX6 U2887 ( .A(n948), .B(n542), .C(n2710), .Z(n2719) );
  AO7CSVTX6 U2888 ( .A(n760), .B(n2728), .C(n1642), .Z(n2142) );
  ND2ASVTX8 U2889 ( .A(n2947), .B(n3014), .Z(n2728) );
  ND2SVTX8 U2890 ( .A(n762), .B(n761), .Z(n4106) );
  AN2SVTX8 U2891 ( .A(n765), .B(n3686), .Z(n1953) );
  ND4SVTX6 U2892 ( .A(n1559), .B(n4136), .C(n3018), .D(n767), .Z(n1075) );
  AO7SVTX8 U2893 ( .A(n3371), .B(n2437), .C(n3334), .Z(n4157) );
  ND3SVTX8 U2894 ( .A(n1982), .B(n482), .C(n3392), .Z(n3334) );
  ND2SVTX8 U2895 ( .A(n1396), .B(n768), .Z(n3371) );
  ND2SVTX6 U2896 ( .A(n3390), .B(n1394), .Z(n768) );
  NR2ASVTX6 U2897 ( .A(n770), .B(n4157), .Z(n769) );
  ND2SVTX4 U2898 ( .A(n3312), .B(n3246), .Z(n4158) );
  NR2SVTX4 U2899 ( .A(n3212), .B(n771), .Z(n2775) );
  ND2SVTX4 U2900 ( .A(n3212), .B(n771), .Z(n3352) );
  AO5ASVTX8 U2901 ( .B(n507), .A(n2774), .C(n2772), .Z(n2801) );
  AO7SVTX6 U2902 ( .A(n402), .B(n1728), .C(n956), .Z(n2771) );
  ND2SVTX4 U2903 ( .A(n772), .B(n2037), .Z(n956) );
  CTIVSVTX4 U2904 ( .A(n774), .Z(n3039) );
  ENSVTX8 U2905 ( .A(n779), .B(n615), .Z(n774) );
  EN3SVTX8 U2906 ( .A(n342), .B(n1764), .C(n1743), .Z(n3005) );
  EO3SVTX8 U2907 ( .A(n1346), .B(n2944), .C(n2945), .Z(n2786) );
  IVSVTX4 U2908 ( .A(n2398), .Z(n777) );
  ND2SVTX6 U2909 ( .A(n780), .B(n2801), .Z(n3337) );
  IVSVTX4 U2910 ( .A(n3726), .Z(n781) );
  ND2ASVTX8 U2911 ( .A(n1352), .B(n556), .Z(n4274) );
  IVSVTX4 U2912 ( .A(n1357), .Z(n1431) );
  AO7SVTX6 U2913 ( .A(n4077), .B(n784), .C(n782), .Z(n1357) );
  ND2SVTX4 U2914 ( .A(n783), .B(n1356), .Z(n782) );
  NR2SVTX4 U2915 ( .A(n3158), .B(n3149), .Z(n783) );
  IVSVTX4 U2916 ( .A(n785), .Z(n3975) );
  ND2ASVTX8 U2917 ( .A(n2381), .B(n3327), .Z(n3376) );
  AO6SVTX2 U2918 ( .A(n792), .B(n791), .C(n4138), .Z(n790) );
  IVSVTX12 U2919 ( .A(n4106), .Z(n2352) );
  ND2SVTX4 U2920 ( .A(n514), .B(n793), .Z(n1630) );
  ND2SVTX4 U2921 ( .A(n794), .B(n832), .Z(n812) );
  AO7SVTX8 U2922 ( .A(n4262), .B(n4261), .C(n797), .Z(n4260) );
  EO3SVTX8 U2923 ( .A(n1121), .B(n519), .C(n625), .Z(n800) );
  AO7SVTX8 U2924 ( .A(n2078), .B(n801), .C(n881), .Z(n907) );
  AO7SVTX8 U2925 ( .A(n3557), .B(n807), .C(n1661), .Z(n3465) );
  BFSVTX12 U2926 ( .A(n807), .Z(n805) );
  AO7SVTX6 U2927 ( .A(n805), .B(n3475), .C(n806), .Z(n1427) );
  ND2SVTX4 U2928 ( .A(n616), .B(n618), .Z(n874) );
  ND3SVTX6 U2929 ( .A(n616), .B(n618), .C(n948), .Z(n2712) );
  ND2SVTX8 U2930 ( .A(n2730), .B(n2729), .Z(n1748) );
  ND2SVTX4 U2931 ( .A(n867), .B(n809), .Z(n828) );
  ND2SVTX4 U2932 ( .A(n3661), .B(n3662), .Z(n810) );
  ND2SVTX4 U2933 ( .A(n3703), .B(n3706), .Z(n811) );
  IVSVTX4 U2934 ( .A(n3703), .Z(n2894) );
  IVSVTX12 U2935 ( .A(n808), .Z(n814) );
  IVSVTX4 U2936 ( .A(n1552), .Z(n840) );
  ND2SVTX4 U2937 ( .A(n2887), .B(n816), .Z(n815) );
  IVSVTX4 U2938 ( .A(n818), .Z(n1102) );
  ND3ASVTX8 U2939 ( .A(n584), .B(n2018), .C(n2981), .Z(n819) );
  NR2SVTX8 U2940 ( .A(n1784), .B(n819), .Z(n2140) );
  ND2SVTX6 U2941 ( .A(n820), .B(n2680), .Z(n1120) );
  EO3SVTX8 U2942 ( .A(n822), .B(n1939), .C(n612), .Z(n2996) );
  ND2SVTX4 U2943 ( .A(n826), .B(n825), .Z(n2419) );
  AO7SVTX6 U2944 ( .A(n823), .B(n691), .C(n3078), .Z(n825) );
  ND2SVTX4 U2945 ( .A(n823), .B(n691), .Z(n826) );
  AO4SVTX8 U2946 ( .A(n827), .B(n1297), .C(n2115), .D(n1872), .Z(n1541) );
  IVSVTX6 U2947 ( .A(n827), .Z(n2676) );
  NR3ABSVTX6 U2948 ( .A(n1081), .B(n3904), .C(n828), .Z(n4215) );
  ND2SVTX8 U2949 ( .A(n1706), .B(n829), .Z(n4216) );
  EO3SVTX8 U2950 ( .A(n609), .B(n2818), .C(n2817), .Z(n833) );
  ND3SVTX8 U2951 ( .A(n2656), .B(n834), .C(n1965), .Z(n2736) );
  AO4SVTX8 U2952 ( .A(n2334), .B(n2902), .C(n2753), .D(n918), .Z(n873) );
  AO6SVTX8 U2953 ( .A(n632), .B(n1287), .C(n835), .Z(n1967) );
  AO5SVTX4 U2954 ( .A(n1967), .B(n2887), .C(n628), .Z(n2858) );
  IVSVTX4 U2955 ( .A(n838), .Z(n3349) );
  ND3SVTX6 U2956 ( .A(n3320), .B(n1401), .C(n1400), .Z(n838) );
  EN3SVTX8 U2957 ( .A(n1268), .B(n1647), .C(n969), .Z(n841) );
  ND2SVTX4 U2958 ( .A(n2456), .B(n3204), .Z(n1317) );
  F_ENSVTX2 U2959 ( .A(n842), .B(n3499), .Z(n3500) );
  ND2SVTX4 U2960 ( .A(n3588), .B(n3594), .Z(n842) );
  IVSVTX4 U2961 ( .A(n3654), .Z(n843) );
  NR2ASVTX6 U2962 ( .A(n565), .B(n2234), .Z(n2277) );
  IVSVTX4 U2963 ( .A(n2737), .Z(n1889) );
  IVSVTX12 U2964 ( .A(n1061), .Z(n1538) );
  AO7SVTX8 U2965 ( .A(n2420), .B(n845), .C(n3525), .Z(n2196) );
  NR2SVTX4 U2966 ( .A(n1087), .B(n3442), .Z(n845) );
  AO17SVTX8 U2967 ( .A(n2117), .B(n4266), .C(n1875), .D(n1874), .Z(n4261) );
  ND2SVTX4 U2968 ( .A(n846), .B(n2645), .Z(n1762) );
  ENSVTX8 U2969 ( .A(n2831), .B(n2068), .Z(n2069) );
  AO7SVTX6 U2970 ( .A(n3049), .B(n1686), .C(n3098), .Z(n3050) );
  ND2SVTX4 U2971 ( .A(n4022), .B(n3845), .Z(n2359) );
  AO4SVTX8 U2972 ( .A(n1767), .B(n2582), .C(n551), .D(n2561), .Z(n1772) );
  ND3SVTX8 U2973 ( .A(n2486), .B(n2577), .C(n2489), .Z(n847) );
  AO7ABSVTX6 U2974 ( .A(n1149), .B(n962), .C(n2850), .Z(n2851) );
  ND4ABSVTX8 U2975 ( .A(n2678), .B(n1231), .C(n2155), .D(n1229), .Z(n2810) );
  ND2ASVTX1 U2976 ( .A(n2512), .B(n2308), .Z(n1564) );
  IVSVTX4 U2977 ( .A(n2266), .Z(n1514) );
  ND3ABSVTX8 U2978 ( .A(n512), .B(n1023), .C(n2180), .Z(n1724) );
  ND2SVTX4 U2979 ( .A(n850), .B(n849), .Z(n2998) );
  ND2SVTX4 U2980 ( .A(n2993), .B(n3283), .Z(n850) );
  EN3SVTX8 U2981 ( .A(n2353), .B(n2993), .C(n851), .Z(n3000) );
  IVSVTX4 U2982 ( .A(n3283), .Z(n851) );
  NR2SVTX4 U2983 ( .A(n854), .B(n853), .Z(n852) );
  NR2SVTX4 U2984 ( .A(n2107), .B(n1696), .Z(n853) );
  ND2SVTX4 U2985 ( .A(n2076), .B(n2108), .Z(n854) );
  AO6ASVTX8 U2986 ( .A(n1297), .B(n2677), .C(n1124), .Z(n1974) );
  AO4SVTX4 U2987 ( .A(n1466), .B(n3513), .C(n2291), .D(n3500), .Z(n1947) );
  IVSVTX4 U2988 ( .A(n2710), .Z(n2309) );
  CTIVSVTX4 U2989 ( .A(n3486), .Z(n1747) );
  IVSVTX12 U2990 ( .A(n3282), .Z(n3068) );
  ND2SVTX8 U2991 ( .A(n2563), .B(n2184), .Z(n2183) );
  ND3SVTX8 U2992 ( .A(n1280), .B(n1284), .C(n1277), .Z(n4086) );
  IVSVTX4 U2993 ( .A(n1164), .Z(n860) );
  IVSVTX12 U2994 ( .A(n1107), .Z(n1023) );
  ND2SVTX4 U2995 ( .A(n555), .B(n1043), .Z(n2674) );
  IVSVTX8 U2996 ( .A(n2514), .Z(n2377) );
  ND2SVTX6 U2997 ( .A(n1540), .B(n1113), .Z(n1539) );
  ND3ASVTX8 U2998 ( .A(n1107), .B(n2630), .C(n1060), .Z(n1916) );
  F_EOSVTX2 U2999 ( .A(n1266), .B(n1690), .Z(n1377) );
  NR3ASVTX8 U3000 ( .A(n878), .B(n2424), .C(n1777), .Z(n4050) );
  ND2SVTX4 U3001 ( .A(n514), .B(n2268), .Z(n864) );
  AO3SVTX6 U3002 ( .A(n1824), .B(n1509), .C(n1510), .D(n4138), .Z(n866) );
  AO7ABSVTX8 U3003 ( .A(n428), .B(n1089), .C(n1815), .Z(n2880) );
  IVSVTX4 U3004 ( .A(n1112), .Z(n1113) );
  EN3SVTX6 U3005 ( .A(n2789), .B(n942), .C(n622), .Z(n2778) );
  IVSVTX4 U3006 ( .A(n3526), .Z(n872) );
  AN2SVTX8 U3007 ( .A(n3525), .B(n872), .Z(n3527) );
  AO2SVTX6 U3008 ( .A(n1377), .B(n561), .C(n1375), .D(n1976), .Z(n1374) );
  IVSVTX12 U3009 ( .A(n873), .Z(n1939) );
  ND2SVTX4 U3010 ( .A(n2802), .B(n2803), .Z(n3382) );
  ND3SVTX8 U3011 ( .A(n955), .B(n3588), .C(n3589), .Z(n1810) );
  IVSVTX4 U3012 ( .A(n2525), .Z(n2298) );
  NR2SVTX4 U3013 ( .A(n963), .B(n2525), .Z(n2226) );
  IVSVTX12 U3014 ( .A(n3273), .Z(n944) );
  ND2SVTX4 U3015 ( .A(n1576), .B(n2899), .Z(n2604) );
  ND2SVTX6 U3016 ( .A(n2819), .B(n2170), .Z(n1798) );
  ND4SVTX4 U3017 ( .A(n3024), .B(n2724), .C(n2725), .D(n598), .Z(n896) );
  IVSVTX4 U3018 ( .A(n3094), .Z(n1236) );
  EN3SVTX8 U3019 ( .A(n611), .B(n609), .C(n506), .Z(n2216) );
  ND2ASVTX8 U3020 ( .A(n2505), .B(n2506), .Z(n1039) );
  IVSVTX2 U3021 ( .A(n3839), .Z(n1305) );
  ND2SVTX4 U3022 ( .A(n2424), .B(n3847), .Z(n2337) );
  ND2SVTX4 U3023 ( .A(n3840), .B(n2120), .Z(n3847) );
  ND3SVTX8 U3024 ( .A(n1378), .B(n1374), .C(n1380), .Z(n954) );
  AO7SVTX6 U3025 ( .A(n3757), .B(n3758), .C(n1683), .Z(n3759) );
  BFSVTX4 U3026 ( .A(n1872), .Z(rslt_o[28]) );
  IVSVTX8 U3027 ( .A(n1269), .Z(n1270) );
  IVSVTX10 U3028 ( .A(n1732), .Z(n2398) );
  IVSVTX4 U3029 ( .A(n2655), .Z(n1761) );
  ND3SVTX8 U3030 ( .A(n622), .B(n1482), .C(n598), .Z(n2088) );
  IVSVTX6 U3031 ( .A(n3865), .Z(n3779) );
  EO3SVTX8 U3032 ( .A(n507), .B(n2773), .C(n2772), .Z(n2803) );
  EOSVTX8 U3033 ( .A(n456), .B(n2850), .Z(n2861) );
  NR2ASVTX6 U3034 ( .A(n3873), .B(n877), .Z(n3875) );
  AO1SVTX8 U3035 ( .A(n2105), .B(n1838), .C(n3794), .D(n494), .Z(n2104) );
  IVSVTX4 U3036 ( .A(n2994), .Z(n1807) );
  NR2SVTX6 U3037 ( .A(n1871), .B(n1765), .Z(n2859) );
  ND2SVTX6 U3038 ( .A(n1584), .B(n1583), .Z(n1106) );
  ND3ABSVTX8 U3039 ( .A(n1939), .B(n1142), .C(n3280), .Z(n2642) );
  CTBUFSVTX4 U3040 ( .A(n343), .Z(n2698) );
  ND2SVTX6 U3041 ( .A(n1937), .B(n3079), .Z(n2147) );
  NR2SVTX4 U3042 ( .A(n728), .B(n2240), .Z(n879) );
  IVSVTX8 U3043 ( .A(n2497), .Z(n2514) );
  BFSVTX8 U3044 ( .A(n2353), .Z(n1669) );
  IVSVTX8 U3045 ( .A(n2812), .Z(n2370) );
  AO17SVTX8 U3046 ( .A(n1684), .B(n1222), .C(n3893), .D(n3885), .Z(n3857) );
  AO4SVTX8 U3047 ( .A(n1544), .B(n1542), .C(n2671), .D(n2294), .Z(n2115) );
  IVSVTX4 U3048 ( .A(n882), .Z(n2012) );
  IVSVTX2 U3049 ( .A(n2787), .Z(n1679) );
  CTIVSVTX4 U3050 ( .A(n2067), .Z(n2233) );
  ND2SVTX4 U3051 ( .A(n793), .B(n3146), .Z(n3163) );
  AO7NSVTX4 U3052 ( .A(n4031), .B(n3401), .C(n3613), .Z(n2408) );
  ND2SVTX4 U3053 ( .A(n3912), .B(n3920), .Z(n3728) );
  NR2SVTX4 U3054 ( .A(n2266), .B(n2323), .Z(n884) );
  ND2SVTX4 U3055 ( .A(n1934), .B(n2108), .Z(n2075) );
  ND2SVTX4 U3056 ( .A(n1648), .B(n886), .Z(n2289) );
  ND2SVTX4 U3057 ( .A(n3964), .B(n974), .Z(n3961) );
  EO3SVTX8 U3058 ( .A(n643), .B(n627), .C(n1937), .Z(n2876) );
  NR2SVTX4 U3059 ( .A(n3106), .B(n525), .Z(n888) );
  AO17SVTX2 U3060 ( .A(n831), .B(n869), .C(n2431), .D(n3689), .Z(n3700) );
  ND4SVTX6 U3061 ( .A(n3721), .B(n3727), .C(n3735), .D(n3736), .Z(n3762) );
  ND3SVTX8 U3062 ( .A(n2561), .B(n2698), .C(n1197), .Z(n2562) );
  ND2SVTX4 U3063 ( .A(n1162), .B(n890), .Z(n894) );
  ND2SVTX4 U3064 ( .A(n563), .B(n1245), .Z(n890) );
  ND4ASVTX8 U3065 ( .A(n606), .B(n3017), .C(n3015), .D(n3016), .Z(n1073) );
  AN2SVTX4 U3066 ( .A(n3817), .B(n3818), .Z(n3872) );
  IVSVTX4 U3067 ( .A(n894), .Z(n1071) );
  AO7SVTX8 U3068 ( .A(n4114), .B(n4113), .C(n4112), .Z(n4206) );
  AO7CSVTX8 U3069 ( .A(n532), .B(n1270), .C(n3140), .Z(n1255) );
  BFSVTX6 U3070 ( .A(n620), .Z(n2129) );
  AO7ABSVTX8 U3071 ( .A(n1233), .B(n1797), .C(n1230), .Z(n2565) );
  ND2ASVTX8 U3072 ( .A(n4101), .B(n1244), .Z(n4141) );
  F_ENSVTX2 U3073 ( .A(n2789), .B(n617), .Z(n1242) );
  NR2SVTX8 U3074 ( .A(n3760), .B(n3759), .Z(n3908) );
  AO7SVTX2 U3075 ( .A(n3551), .B(n2419), .C(n3550), .Z(n3556) );
  ND3SVTX8 U3076 ( .A(n3522), .B(n2763), .C(n2987), .Z(n3594) );
  AO4SVTX8 U3077 ( .A(n2704), .B(n1287), .C(n2902), .D(n2143), .Z(n2255) );
  ND2SVTX4 U3078 ( .A(n1083), .B(n2806), .Z(n1527) );
  ND2SVTX4 U3079 ( .A(n1049), .B(n2831), .Z(n2832) );
  AO20SVTX8 U3080 ( .A(n898), .B(n3349), .C(n3382), .D(n1097), .Z(n978) );
  AO2ASVTX6 U3081 ( .C(n2661), .D(n1336), .A(n1107), .B(n1233), .Z(n966) );
  ND2ASVTX8 U3082 ( .A(n3529), .B(n1876), .Z(n4266) );
  ND2SVTX6 U3083 ( .A(n3907), .B(n3906), .Z(n4213) );
  EO3SVTX8 U3084 ( .A(n520), .B(n2843), .C(n2842), .Z(n3483) );
  AO20SVTX8 U3085 ( .A(n1158), .B(n1157), .C(n4136), .D(n2828), .Z(n1074) );
  F_EOSVTX2 U3086 ( .A(n4014), .B(n3604), .Z(n3605) );
  BFSVTX1 U3087 ( .A(n1219), .Z(rslt_o[30]) );
  AO7ABSVTX8 U3088 ( .A(n728), .B(n1438), .C(n2842), .Z(n1437) );
  ND2SVTX4 U3089 ( .A(n903), .B(n2687), .Z(n902) );
  ND3SVTX8 U3090 ( .A(n2118), .B(n1322), .C(n1082), .Z(n2368) );
  NR2SVTX4 U3091 ( .A(n3887), .B(n3832), .Z(n906) );
  IVSVTX10 U3092 ( .A(n4106), .Z(n1777) );
  AO7ABSVTX4 U3093 ( .A(n1608), .B(n1609), .C(n2748), .Z(n2757) );
  IVSVTX4 U3094 ( .A(n1263), .Z(n1262) );
  F_EOSVTX2 U3095 ( .A(n1346), .B(n1347), .Z(n1348) );
  ND3ABSVTX8 U3096 ( .A(n3903), .B(n586), .C(n3948), .Z(n908) );
  ND4SVTX4 U3097 ( .A(n3903), .B(n4022), .C(n1970), .D(n3845), .Z(n909) );
  ND2SVTX2 U3098 ( .A(n2534), .B(n2126), .Z(n2535) );
  IVSVTX4 U3099 ( .A(n3251), .Z(n910) );
  EO3SVTX8 U3100 ( .A(n2849), .B(n627), .C(n1472), .Z(n2850) );
  AO6SVTX4 U3101 ( .A(n912), .B(num_i[3]), .C(n2510), .Z(n2511) );
  BFSVTX2 U3102 ( .A(n4291), .Z(n1731) );
  IVSVTX6 U3103 ( .A(n2014), .Z(n4022) );
  ND2ASVTX8 U3104 ( .A(n2014), .B(n3845), .Z(n2239) );
  ND2SVTX4 U3105 ( .A(n913), .B(n2521), .Z(n2544) );
  BFSVTX8 U3106 ( .A(n1025), .Z(n1030) );
  IVSVTX4 U3107 ( .A(num_i[17]), .Z(n1941) );
  ND2SVTX4 U3108 ( .A(n2578), .B(n892), .Z(n2520) );
  AO7SVTX4 U3109 ( .A(n709), .B(n1372), .C(n1647), .Z(n2840) );
  NR2ASVTX6 U3110 ( .A(n1978), .B(n2914), .Z(n1977) );
  ND3ASVTX6 U3111 ( .A(n555), .B(n1047), .C(n1026), .Z(n2760) );
  F_ENSVTX2 U3112 ( .A(n3497), .B(n3496), .Z(n1627) );
  ND4ABSVTX8 U3113 ( .A(n865), .B(n916), .C(n496), .D(n1467), .Z(n1775) );
  ND2SVTX4 U3114 ( .A(n917), .B(n2623), .Z(n2567) );
  NR2SVTX4 U3115 ( .A(n1107), .B(n1538), .Z(n917) );
  NR4ABCSVTX6 U3116 ( .A(n1361), .B(n502), .C(n608), .D(n610), .Z(n2738) );
  ND2SVTX4 U3117 ( .A(n549), .B(n2110), .Z(n2593) );
  ND2ASVTX8 U3118 ( .A(n919), .B(n2146), .Z(n2994) );
  AO2SVTX8 U3119 ( .A(n2610), .B(n950), .C(n2403), .D(n1894), .Z(n2560) );
  AO3SVTX8 U3120 ( .A(rslt_o[31]), .B(n2537), .C(n2535), .D(n2536), .Z(n2610)
         );
  EN3SVTX8 U3121 ( .A(n1669), .B(n620), .C(n962), .Z(n3094) );
  ND2SVTX4 U3122 ( .A(n921), .B(n1640), .Z(n3614) );
  IVSVTX4 U3123 ( .A(n3445), .Z(n1123) );
  NR2SVTX4 U3124 ( .A(n3810), .B(n928), .Z(n3632) );
  ND2SVTX4 U3125 ( .A(n4031), .B(n3401), .Z(n3399) );
  IVSVTX6 U3126 ( .A(n1319), .Z(n3391) );
  ND2ASVTX8 U3127 ( .A(n3122), .B(n3055), .Z(n3393) );
  NR2SVTX6 U3128 ( .A(n1716), .B(n931), .Z(n1391) );
  ENSVTX8 U3129 ( .A(n941), .B(n3046), .Z(n3396) );
  IVSVTX4 U3130 ( .A(n942), .Z(n1892) );
  NR2SVTX8 U3131 ( .A(n1481), .B(n943), .Z(n2664) );
  EN3SVTX8 U3132 ( .A(n519), .B(n943), .C(n541), .Z(n993) );
  EN3SVTX8 U3133 ( .A(n943), .B(n1143), .C(n1764), .Z(n959) );
  NR2SVTX8 U3134 ( .A(n1022), .B(n1996), .Z(n951) );
  AO5SVTX4 U3135 ( .A(n1526), .B(n948), .C(n617), .Z(n1334) );
  ND3SVTX8 U3136 ( .A(n955), .B(n3591), .C(n3590), .Z(n3592) );
  ND2ASVTX8 U3137 ( .A(n2994), .B(n2992), .Z(n955) );
  ENSVTX8 U3138 ( .A(n1005), .B(n956), .Z(n2805) );
  ND2SVTX4 U3139 ( .A(n1173), .B(n957), .Z(n2222) );
  ND2ASVTX8 U3140 ( .A(n536), .B(n3998), .Z(n1173) );
  ND3SVTX6 U3141 ( .A(n552), .B(n1805), .C(n1061), .Z(n2665) );
  EN3SVTX8 U3142 ( .A(n728), .B(n2822), .C(n993), .Z(n3839) );
  AO17ASVTX8 U3143 ( .A(n3282), .B(n996), .C(n959), .D(n995), .Z(n2829) );
  AO7ABSVTX8 U3144 ( .A(n1529), .B(n501), .C(n1537), .Z(n2822) );
  AO5ASVTX8 U3145 ( .B(n1664), .A(n520), .C(n958), .Z(n2821) );
  NR2SVTX8 U3146 ( .A(n463), .B(n994), .Z(n997) );
  ND2SVTX8 U3147 ( .A(n3003), .B(n3002), .Z(n961) );
  ND3ABSVTX8 U3148 ( .A(n1635), .B(n1316), .C(n961), .Z(n3015) );
  ND2SVTX4 U3149 ( .A(n567), .B(n961), .Z(n4122) );
  ND2SVTX4 U3150 ( .A(n814), .B(n962), .Z(n2969) );
  ND2SVTX4 U3151 ( .A(n962), .B(n2855), .Z(n2856) );
  ND2SVTX8 U3152 ( .A(n2193), .B(n2192), .Z(n963) );
  AO2SVTX8 U3153 ( .A(n968), .B(n967), .C(n2677), .D(n1323), .Z(n2639) );
  AO2ABSVTX8 U3154 ( .C(n2635), .D(n2634), .A(n2294), .B(n554), .Z(n2677) );
  IVSVTX12 U3155 ( .A(n972), .Z(n1061) );
  ND3SVTX8 U3156 ( .A(n973), .B(n2320), .C(n1092), .Z(n972) );
  NR2SVTX8 U3157 ( .A(n2485), .B(n2484), .Z(n2320) );
  ND3SVTX8 U3158 ( .A(n2477), .B(n2531), .C(n2476), .Z(n1092) );
  NR2SVTX8 U3159 ( .A(n3959), .B(n3957), .Z(n3866) );
  ND4ABCSVTX8 U3160 ( .A(n1785), .B(n3866), .C(n3779), .D(n2374), .Z(n2981) );
  ND2ASVTX8 U3161 ( .A(n1711), .B(n2976), .Z(n2374) );
  ND2SVTX4 U3162 ( .A(n2190), .B(n2020), .Z(n2018) );
  NR2SVTX6 U3163 ( .A(num_i[8]), .B(num_i[9]), .Z(n2193) );
  ND2SVTX4 U3164 ( .A(n3364), .B(n2272), .Z(n976) );
  IVSVTX4 U3165 ( .A(n984), .Z(n977) );
  AO1SVTX6 U3166 ( .A(n489), .B(n980), .C(n979), .D(n978), .Z(n983) );
  NR2SVTX4 U3167 ( .A(n1097), .B(n984), .Z(n980) );
  IVSVTX4 U3168 ( .A(n2135), .Z(n984) );
  IVSVTX4 U3169 ( .A(n1920), .Z(n986) );
  ND2SVTX8 U3170 ( .A(n988), .B(n1179), .Z(n1178) );
  ND3SVTX8 U3171 ( .A(n988), .B(n1179), .C(n2678), .Z(n2679) );
  ND2SVTX8 U3172 ( .A(n3956), .B(n3722), .Z(n3977) );
  ND4SVTX8 U3173 ( .A(n2545), .B(n2547), .C(n992), .D(n1701), .Z(n2532) );
  ND2SVTX8 U3174 ( .A(n1936), .B(n2308), .Z(n992) );
  ND2SVTX6 U3175 ( .A(n998), .B(n999), .Z(n1048) );
  AO6SVTX6 U3176 ( .A(n2576), .B(n2548), .C(n1001), .Z(n1000) );
  NR2ASVTX6 U3177 ( .A(n2348), .B(n3310), .Z(n3048) );
  IVSVTX12 U3178 ( .A(n1002), .Z(n1090) );
  ND2SVTX8 U3179 ( .A(n2680), .B(n1026), .Z(n2729) );
  ND2SVTX8 U3180 ( .A(n2982), .B(n2279), .Z(n2730) );
  AO7SVTX6 U3181 ( .A(n1651), .B(n2306), .C(n1995), .Z(n1003) );
  ENSVTX8 U3182 ( .A(n2805), .B(n1007), .Z(n3998) );
  ND2SVTX4 U3183 ( .A(n1173), .B(n3999), .Z(n4021) );
  AO7SVTX6 U3184 ( .A(n478), .B(n2185), .C(n1416), .Z(n1004) );
  ENSVTX8 U3185 ( .A(n1346), .B(n1006), .Z(n1005) );
  F_ENSVTX2 U3186 ( .A(n3111), .B(n2348), .Z(n1007) );
  ND2SVTX4 U3187 ( .A(n4025), .B(n2430), .Z(n1012) );
  ND2ASVTX8 U3188 ( .A(n4051), .B(n1582), .Z(n4278) );
  ND4ABSVTX8 U3189 ( .A(n1184), .B(n1183), .C(n1189), .D(n1188), .Z(n1582) );
  ND2SVTX6 U3190 ( .A(n4219), .B(n1008), .Z(n4052) );
  ND4SVTX6 U3191 ( .A(n583), .B(n4003), .C(n2135), .D(n4002), .Z(n1013) );
  ND2SVTX4 U3192 ( .A(n1013), .B(n1673), .Z(n1010) );
  ND2SVTX4 U3193 ( .A(n2364), .B(n1015), .Z(n2635) );
  ND2SVTX8 U3194 ( .A(n1586), .B(n1585), .Z(n1015) );
  ND2SVTX6 U3195 ( .A(n2120), .B(n1018), .Z(n1017) );
  NR2SVTX6 U3196 ( .A(n2829), .B(n3839), .Z(n1018) );
  ND4SVTX8 U3197 ( .A(n1137), .B(n1141), .C(n1139), .D(n1136), .Z(n1020) );
  IVSVTX4 U3198 ( .A(n1020), .Z(n3560) );
  ND2ASVTX8 U3199 ( .A(n522), .B(n1020), .Z(n4257) );
  ND2SVTX6 U3200 ( .A(n1023), .B(n1061), .Z(n1421) );
  AO7ABSVTX8 U3201 ( .A(n1762), .B(n1872), .C(n1167), .Z(n2982) );
  ND2SVTX8 U3202 ( .A(n2730), .B(n2729), .Z(n1025) );
  NR2SVTX4 U3203 ( .A(n1029), .B(n1027), .Z(n1190) );
  AO6SVTX4 U3204 ( .A(n1530), .B(n3996), .C(n3946), .Z(n1029) );
  ND2SVTX8 U3205 ( .A(n1032), .B(n1031), .Z(n1388) );
  NR2SVTX8 U3206 ( .A(num_i[12]), .B(num_i[15]), .Z(n1032) );
  ND2SVTX6 U3207 ( .A(n3504), .B(n3503), .Z(n1128) );
  ND2SVTX4 U3208 ( .A(n1580), .B(n1034), .Z(n2592) );
  ND2SVTX6 U3209 ( .A(n2609), .B(n950), .Z(n2602) );
  AO2SVTX6 U3210 ( .A(n2289), .B(n950), .C(n418), .D(n2700), .Z(n2307) );
  NR2SVTX4 U3211 ( .A(n638), .B(n1768), .Z(n1037) );
  ND2SVTX4 U3212 ( .A(n2504), .B(n1038), .Z(n2505) );
  IVSVTX4 U3213 ( .A(n2722), .Z(n2721) );
  ND2ASVTX8 U3214 ( .A(n2880), .B(n1041), .Z(n3706) );
  ND2SVTX6 U3215 ( .A(n1521), .B(n3070), .Z(n1661) );
  ND2ASVTX8 U3216 ( .A(n1522), .B(n3066), .Z(n1521) );
  IVSVTX4 U3217 ( .A(n1661), .Z(n3461) );
  ND2SVTX4 U3218 ( .A(n2643), .B(n2070), .Z(n1045) );
  AO17SVTX6 U3219 ( .A(n1715), .B(n1562), .C(n1075), .D(n1046), .Z(n1069) );
  NR2SVTX8 U3220 ( .A(n1074), .B(n1070), .Z(n1046) );
  ND2SVTX4 U3221 ( .A(n2900), .B(n1048), .Z(n3271) );
  AO7SVTX6 U3222 ( .A(n1360), .B(n2666), .C(n2665), .Z(n2753) );
  ND2SVTX4 U3223 ( .A(n472), .B(n1052), .Z(n1051) );
  ND2SVTX4 U3224 ( .A(n1053), .B(n2959), .Z(n3323) );
  IVSVTX4 U3225 ( .A(n2960), .Z(n1053) );
  ND2SVTX6 U3226 ( .A(n2957), .B(n2958), .Z(n2962) );
  EN3SVTX6 U3227 ( .A(n518), .B(n617), .C(n2868), .Z(n2963) );
  AO2SVTX8 U3228 ( .A(n2703), .B(n2902), .C(n2705), .D(n2576), .Z(n1642) );
  ND4SVTX8 U3229 ( .A(n1055), .B(n1057), .C(n1054), .D(n1056), .Z(n2705) );
  ND2SVTX6 U3230 ( .A(n2587), .B(n2681), .Z(n1054) );
  AO7ABSVTX8 U3231 ( .A(rslt_o[28]), .B(n2048), .C(n1534), .Z(n2703) );
  ND2SVTX4 U3232 ( .A(n1580), .B(n2036), .Z(n1057) );
  IVSVTX4 U3233 ( .A(n1059), .Z(n2833) );
  ND2SVTX8 U3234 ( .A(n2679), .B(n1200), .Z(n1199) );
  AO3SVTX6 U3235 ( .A(n1062), .B(n2892), .C(n1794), .D(n2891), .Z(n3663) );
  AO1CDSVTX8 U3236 ( .A(n3663), .B(n1063), .C(n3706), .D(n3703), .Z(n3415) );
  NR2ASVTX6 U3237 ( .A(n2891), .B(n613), .Z(n3487) );
  AO7SVTX8 U3238 ( .A(n1986), .B(n1064), .C(n3573), .Z(n1489) );
  IVSVTX4 U3239 ( .A(n2649), .Z(n1067) );
  ND4ABSVTX8 U3240 ( .A(n1067), .B(n2678), .C(n2650), .D(n2648), .Z(n2735) );
  IVSVTX2 U3241 ( .A(n3724), .Z(n3004) );
  ND2ASVTX8 U3242 ( .A(n3007), .B(n3008), .Z(n3420) );
  NR2SVTX8 U3243 ( .A(n600), .B(n1078), .Z(n3422) );
  AO7SVTX6 U3244 ( .A(n3006), .B(n3005), .C(n3724), .Z(n1078) );
  AO6ASVTX8 U3245 ( .A(n1488), .B(n3420), .C(n1077), .Z(n2442) );
  NR3SVTX8 U3246 ( .A(n3907), .B(n3868), .C(n3869), .Z(n1082) );
  AO2SVTX6 U3247 ( .A(n2239), .B(n462), .C(n3825), .D(n3826), .Z(n2118) );
  ND3ABSVTX8 U3248 ( .A(n2631), .B(n1769), .C(n2636), .Z(n2666) );
  BFSVTX10 U3249 ( .A(n900), .Z(n1083) );
  IVSVTX4 U3250 ( .A(n2334), .Z(n2838) );
  IVSVTX4 U3251 ( .A(n2678), .Z(n2839) );
  ND2SVTX4 U3252 ( .A(n684), .B(n2352), .Z(n2748) );
  NR2ASVTX6 U3253 ( .A(n2678), .B(n2565), .Z(n2569) );
  ND2SVTX6 U3254 ( .A(n3442), .B(n1087), .Z(n3525) );
  ND2SVTX8 U3255 ( .A(n3570), .B(n1085), .Z(n3620) );
  F_ENSVTX2 U3256 ( .A(n3572), .B(n1086), .Z(n2268) );
  ND2SVTX4 U3257 ( .A(n3620), .B(n3571), .Z(n1086) );
  IVSVTX4 U3258 ( .A(n2344), .Z(n2387) );
  EN3SVTX8 U3259 ( .A(n619), .B(n1529), .C(n1361), .Z(n2972) );
  NR2SVTX4 U3260 ( .A(n535), .B(n3686), .Z(n3967) );
  ND3ASVTX6 U3261 ( .A(n635), .B(n1904), .C(n2231), .Z(n2594) );
  ND4SVTX4 U3262 ( .A(n2044), .B(n2047), .C(n2175), .D(n2038), .Z(n1351) );
  ND2SVTX6 U3263 ( .A(n1155), .B(n1154), .Z(n2704) );
  ND2SVTX6 U3264 ( .A(n2057), .B(n2407), .Z(n2143) );
  ND2SVTX8 U3265 ( .A(n1252), .B(n1253), .Z(n2784) );
  ND2SVTX1 U3266 ( .A(n4247), .B(n1093), .Z(n4253) );
  IVSVTX4 U3267 ( .A(n2613), .Z(n1094) );
  ND2SVTX4 U3268 ( .A(n2013), .B(n2582), .Z(n1096) );
  ND2SVTX6 U3269 ( .A(n2424), .B(n1111), .Z(n1110) );
  IVSVTX12 U3270 ( .A(n1117), .Z(n1107) );
  ND3SVTX8 U3271 ( .A(n2531), .B(n2226), .C(n2227), .Z(n1108) );
  ENSVTX8 U3272 ( .A(n2420), .B(n3527), .Z(n1111) );
  ND2SVTX2 U3273 ( .A(n1117), .B(n972), .Z(n1118) );
  ND2ASVTX6 U3274 ( .A(n2898), .B(n2183), .Z(n2601) );
  ND2SVTX4 U3275 ( .A(n2590), .B(n2591), .Z(n2598) );
  ND3ABSVTX8 U3276 ( .A(n1861), .B(n2364), .C(n1323), .Z(n2070) );
  IVSVTX4 U3277 ( .A(n3572), .Z(n1122) );
  IVSVTX4 U3278 ( .A(n1986), .Z(n3444) );
  AO3SVTX6 U3279 ( .A(n1123), .B(n1986), .C(n3446), .D(n3573), .Z(n3447) );
  IVSVTX12 U3280 ( .A(n1760), .Z(n1124) );
  ND3SVTX8 U3281 ( .A(n2390), .B(n2012), .C(n471), .Z(n1760) );
  ND3SVTX8 U3282 ( .A(n2474), .B(n2473), .C(n2499), .Z(n2515) );
  ND3SVTX6 U3283 ( .A(n1941), .B(n2577), .C(n2133), .Z(n2516) );
  ND4SVTX4 U3284 ( .A(num_i[11]), .B(n1941), .C(n2577), .D(n2133), .Z(n1125)
         );
  NR2SVTX8 U3285 ( .A(n1388), .B(n2389), .Z(n2531) );
  ND2SVTX6 U3286 ( .A(n2220), .B(n2497), .Z(n2389) );
  ND3ASVTX6 U3287 ( .A(n1125), .B(n2531), .C(n1126), .Z(n2545) );
  ND2SVTX8 U3288 ( .A(n2670), .B(n2669), .Z(n1127) );
  AO7SVTX2 U3289 ( .A(n2459), .B(n3523), .C(n1128), .Z(n3506) );
  ND4SVTX4 U3290 ( .A(n3548), .B(n3549), .C(n3547), .D(n3546), .Z(n1141) );
  ND2ASVTX8 U3291 ( .A(n3531), .B(n745), .Z(n1132) );
  AO21SVTX6 U3292 ( .A(n3620), .B(n3530), .C(n373), .D(n2424), .Z(n1135) );
  ND2SVTX4 U3293 ( .A(n1422), .B(n1138), .Z(n1137) );
  F_ENSVTX2 U3294 ( .A(n2464), .B(n3558), .Z(n1138) );
  AO1CSVTX8 U3295 ( .A(n4066), .B(n3559), .C(n1140), .D(n3537), .Z(n1139) );
  ND2SVTX4 U3296 ( .A(n537), .B(n1710), .Z(n1434) );
  ND2SVTX4 U3297 ( .A(n3704), .B(n1040), .Z(n3664) );
  ND2SVTX4 U3298 ( .A(n543), .B(n2285), .Z(n3062) );
  AO7SVTX6 U3299 ( .A(n1149), .B(n729), .C(n2761), .Z(n2985) );
  AO7SVTX6 U3300 ( .A(n1149), .B(n2970), .C(n2969), .Z(n1771) );
  ND3SVTX6 U3301 ( .A(n2576), .B(n1155), .C(n1154), .Z(n1253) );
  ND2SVTX4 U3302 ( .A(n1156), .B(n2345), .Z(n3020) );
  AO6ASVTX8 U3303 ( .A(n4092), .B(n1557), .C(n2942), .Z(n4136) );
  AO6SVTX4 U3304 ( .A(n3016), .B(n3015), .C(n3014), .Z(n1163) );
  AO7SVTX6 U3305 ( .A(n3014), .B(n3017), .C(n733), .Z(n1164) );
  ND2SVTX4 U3306 ( .A(n4247), .B(n4249), .Z(n3563) );
  ND2SVTX4 U3307 ( .A(n2115), .B(n1538), .Z(n2643) );
  IVSVTX4 U3308 ( .A(n1271), .Z(n1170) );
  ND2SVTX8 U3309 ( .A(n1168), .B(n1169), .Z(n1271) );
  ND2SVTX4 U3310 ( .A(n2923), .B(n1171), .Z(n3301) );
  ND2SVTX4 U3311 ( .A(n2922), .B(n2921), .Z(n3366) );
  ND2ASVTX6 U3312 ( .A(n4149), .B(n1174), .Z(n1659) );
  ND3SVTX8 U3313 ( .A(n4165), .B(n1441), .C(n499), .Z(n1174) );
  ND3SVTX4 U3314 ( .A(n4206), .B(n2421), .C(n1174), .Z(n1599) );
  ND2SVTX4 U3315 ( .A(n1175), .B(n4058), .Z(n1504) );
  ND3ASVTX6 U3316 ( .A(n4143), .B(n1175), .C(n433), .Z(n2005) );
  ND2SVTX8 U3317 ( .A(n2061), .B(n1246), .Z(n4058) );
  ND2SVTX6 U3318 ( .A(n1227), .B(n1997), .Z(n1179) );
  ND2SVTX4 U3319 ( .A(n1187), .B(n1186), .Z(n1185) );
  ND2SVTX4 U3320 ( .A(n3967), .B(n3968), .Z(n1186) );
  NR2SVTX8 U3321 ( .A(num_i[26]), .B(num_i[25]), .Z(n2499) );
  NR2SVTX6 U3322 ( .A(num_i[28]), .B(num_i[24]), .Z(n1198) );
  NR2SVTX8 U3323 ( .A(n4147), .B(n4268), .Z(n1202) );
  ND2SVTX8 U3324 ( .A(n3912), .B(n387), .Z(n3981) );
  ND2SVTX8 U3325 ( .A(n1907), .B(n1906), .Z(n3912) );
  ND2SVTX6 U3326 ( .A(n3411), .B(n3980), .Z(n2920) );
  ND2SVTX8 U3327 ( .A(n599), .B(n2907), .Z(n3980) );
  EN3SVTX6 U3328 ( .A(n948), .B(n618), .C(n1791), .Z(n2339) );
  AO4ABSVTX6 U3329 ( .C(n1728), .D(n2896), .A(n3270), .B(n2017), .Z(n2911) );
  AO7SVTX6 U3330 ( .A(n2971), .B(n1601), .C(n1207), .Z(n1978) );
  NR2SVTX6 U3331 ( .A(n2511), .B(n1209), .Z(n2227) );
  NR2SVTX4 U3332 ( .A(n3686), .B(n1215), .Z(n1214) );
  F_ENSVTX2 U3333 ( .A(n3491), .B(n3490), .Z(n1215) );
  AO7SVTX6 U3334 ( .A(n2077), .B(n3920), .C(n3911), .Z(n3982) );
  ND2SVTX6 U3335 ( .A(n2358), .B(n1884), .Z(n2078) );
  IVSVTX4 U3336 ( .A(n2915), .Z(n1222) );
  ND2SVTX4 U3337 ( .A(n1223), .B(n2807), .Z(n1226) );
  NR2SVTX4 U3338 ( .A(n2660), .B(n512), .Z(n1227) );
  ND2SVTX4 U3339 ( .A(n2636), .B(n2651), .Z(n1228) );
  IVSVTX6 U3340 ( .A(n2565), .Z(n1229) );
  NR2SVTX6 U3341 ( .A(n1421), .B(n1893), .Z(n1231) );
  AO3SVTX8 U3342 ( .A(n2385), .B(n2964), .C(n3323), .D(n3324), .Z(n3206) );
  ENSVTX8 U3343 ( .A(n2954), .B(n2955), .Z(n2964) );
  AO7ABSVTX8 U3344 ( .A(n1932), .B(n615), .C(n1232), .Z(n2954) );
  ND2SVTX8 U3345 ( .A(n2502), .B(n2501), .Z(n1233) );
  ND2SVTX6 U3346 ( .A(n4283), .B(n4305), .Z(n4291) );
  ND2ASVTX8 U3347 ( .A(n2394), .B(n1908), .Z(n4305) );
  NR3SVTX8 U3348 ( .A(n1845), .B(n1841), .C(n1844), .Z(n1234) );
  ND2SVTX4 U3349 ( .A(n3400), .B(n562), .Z(n3406) );
  IVSVTX4 U3350 ( .A(n1238), .Z(n3870) );
  AO7SVTX8 U3351 ( .A(n2573), .B(n2584), .C(n1239), .Z(n2483) );
  AO8SVTX4 U3352 ( .A(n2573), .B(n2518), .C(n2377), .D(n891), .Z(n1675) );
  NR4SVTX6 U3353 ( .A(num_i[11]), .B(num_i[7]), .C(num_i[10]), .D(num_i[6]), 
        .Z(n2470) );
  ND2SVTX8 U3354 ( .A(n2811), .B(n2810), .Z(n2812) );
  IVSVTX4 U3355 ( .A(n1244), .Z(n1243) );
  ND2SVTX4 U3356 ( .A(n2061), .B(n1246), .Z(n1245) );
  ND2SVTX8 U3357 ( .A(n1264), .B(n564), .Z(n2061) );
  ND2SVTX4 U3358 ( .A(n1249), .B(n1248), .Z(n1247) );
  ND2SVTX4 U3359 ( .A(n4306), .B(n4192), .Z(n1248) );
  IVSVTX4 U3360 ( .A(n4272), .Z(n4306) );
  AO6SVTX4 U3361 ( .A(n4289), .B(n1731), .C(n1250), .Z(n1249) );
  IVSVTX4 U3362 ( .A(n540), .Z(n1251) );
  AO7ABSVTX4 U3363 ( .A(n4058), .B(n3309), .C(n1988), .Z(n1987) );
  AO17SVTX4 U3364 ( .A(n2092), .B(n432), .C(n1251), .D(n2164), .Z(n2960) );
  EN3SVTX8 U3365 ( .A(n622), .B(n2945), .C(n624), .Z(n2924) );
  IVSVTX4 U3366 ( .A(n2784), .Z(n1790) );
  ND2SVTX4 U3367 ( .A(n4055), .B(n581), .Z(n1365) );
  ND2SVTX8 U3368 ( .A(n3815), .B(n3814), .Z(n1259) );
  ND2SVTX4 U3369 ( .A(n3171), .B(n1259), .Z(n3172) );
  F_ENSVTX2 U3370 ( .A(n3682), .B(n1863), .Z(n3683) );
  IVSVTX12 U3371 ( .A(n1268), .Z(n3065) );
  ND2SVTX8 U3372 ( .A(n3628), .B(n3629), .Z(n1690) );
  NR2SVTX4 U3373 ( .A(n1278), .B(n1275), .Z(n1277) );
  IVSVTX4 U3374 ( .A(n1279), .Z(n1276) );
  ND4ABSVTX6 U3375 ( .A(n1283), .B(n532), .C(n4058), .D(n4105), .Z(n1282) );
  ND2ASVTX8 U3376 ( .A(n2653), .B(n2256), .Z(n2654) );
  AO17SVTX4 U3377 ( .A(n4059), .B(n1641), .C(n1289), .D(n1290), .Z(n4065) );
  ND2SVTX4 U3378 ( .A(n1289), .B(n4059), .Z(n1290) );
  ND2ASVTX8 U3379 ( .A(n1292), .B(n1705), .Z(n3294) );
  AO7ABSVTX4 U3380 ( .A(n390), .B(n2789), .C(n3038), .Z(n1294) );
  IVSVTX4 U3381 ( .A(n1296), .Z(n3265) );
  NR2SVTX6 U3382 ( .A(n1787), .B(n1296), .Z(n1784) );
  ND2SVTX4 U3383 ( .A(n3265), .B(n3326), .Z(n3327) );
  AO3SVTX6 U3384 ( .A(n3808), .B(n3092), .C(n1299), .D(n3809), .Z(n2204) );
  ND2SVTX8 U3385 ( .A(n3060), .B(n3090), .Z(n1299) );
  IVSVTX4 U3386 ( .A(n1298), .Z(n3631) );
  NR2ASVTX6 U3387 ( .A(n3818), .B(n3874), .Z(n1298) );
  NR2SVTX6 U3388 ( .A(n3247), .B(n1300), .Z(n3178) );
  IVSVTX4 U3389 ( .A(n3244), .Z(n1300) );
  IVSVTX4 U3390 ( .A(n3247), .Z(n3170) );
  ND2SVTX6 U3391 ( .A(n3199), .B(n3198), .Z(n1304) );
  NR3SVTX8 U3392 ( .A(n2195), .B(n1304), .C(n1357), .Z(n1981) );
  ND2ASVTX8 U3393 ( .A(n2829), .B(n1305), .Z(n1499) );
  NR3SVTX8 U3394 ( .A(n1311), .B(n1309), .C(n1306), .Z(n3868) );
  ND2SVTX4 U3395 ( .A(n1313), .B(n1690), .Z(n1308) );
  ND2ASVTX8 U3396 ( .A(n3779), .B(n3960), .Z(n1314) );
  AO7SVTX8 U3397 ( .A(n4119), .B(n531), .C(n3322), .Z(n3204) );
  ND3ABSVTX8 U3398 ( .A(n1315), .B(n509), .C(n3013), .Z(n3016) );
  IVSVTX4 U3399 ( .A(n4175), .Z(n3013) );
  ND3SVTX6 U3400 ( .A(n2456), .B(n1790), .C(n3012), .Z(n1316) );
  ND2ASVTX8 U3401 ( .A(n622), .B(n3143), .Z(n3017) );
  ND3ABSVTX8 U3402 ( .A(n2948), .B(n1318), .C(n1317), .Z(n3143) );
  NR2SVTX4 U3403 ( .A(n2949), .B(n3151), .Z(n1318) );
  NR2SVTX6 U3404 ( .A(n1320), .B(n3056), .Z(n1319) );
  ND2SVTX4 U3405 ( .A(n2092), .B(n2017), .Z(n3044) );
  NR2SVTX4 U3406 ( .A(n2092), .B(n2017), .Z(n3043) );
  AO17DSVTX8 U3407 ( .A(n1023), .B(n2661), .C(n2660), .D(n1061), .Z(n2669) );
  ND2SVTX4 U3408 ( .A(n2829), .B(n3839), .Z(n1325) );
  AO7SVTX8 U3409 ( .A(n1004), .B(n3998), .C(n3927), .Z(n1329) );
  IVSVTX4 U3410 ( .A(n1526), .Z(n1330) );
  IVSVTX4 U3411 ( .A(n1337), .Z(n2428) );
  ND2SVTX4 U3412 ( .A(n583), .B(n3802), .Z(n1337) );
  IVSVTX6 U3413 ( .A(n1341), .Z(n1585) );
  ND3SVTX8 U3414 ( .A(n1479), .B(n1478), .C(n1477), .Z(n1341) );
  ND2ASVTX8 U3415 ( .A(n2825), .B(n1517), .Z(n3927) );
  EO3SVTX8 U3416 ( .A(n1143), .B(n944), .C(n942), .Z(n2817) );
  ND2SVTX4 U3417 ( .A(n567), .B(n3150), .Z(n3153) );
  NR2SVTX6 U3418 ( .A(n4138), .B(n1777), .Z(n3972) );
  EO3SVTX8 U3419 ( .A(n808), .B(n625), .C(n3270), .Z(n1835) );
  ENSVTX4 U3420 ( .A(n1348), .B(n611), .Z(n3011) );
  NR3ABSVTX8 U3421 ( .A(n2044), .B(n2047), .C(n1349), .Z(n1352) );
  NR2ASVTX6 U3422 ( .A(n570), .B(n480), .Z(n2451) );
  ND2ASVTX8 U3423 ( .A(n2975), .B(n2974), .Z(n3626) );
  ND2SVTX6 U3424 ( .A(n2662), .B(n2125), .Z(n1358) );
  ND2SVTX6 U3425 ( .A(n1358), .B(n545), .Z(n2112) );
  IVSVTX12 U3426 ( .A(n2737), .Z(n1361) );
  ND2SVTX8 U3427 ( .A(n2735), .B(n2736), .Z(n2737) );
  ND2SVTX6 U3428 ( .A(n1363), .B(n1362), .Z(n3046) );
  IVSVTX4 U3429 ( .A(n2351), .Z(n2083) );
  NR2SVTX6 U3430 ( .A(n4057), .B(n1365), .Z(n3142) );
  ND2SVTX4 U3431 ( .A(n2911), .B(n1366), .Z(n3412) );
  ND2SVTX4 U3432 ( .A(n2061), .B(n1246), .Z(n2362) );
  ND2ASVTX8 U3433 ( .A(n1368), .B(n1835), .Z(n3093) );
  ND2SVTX8 U3434 ( .A(n1369), .B(n1370), .Z(n3458) );
  AO7ABSVTX8 U3435 ( .A(n401), .B(n3169), .C(n1371), .Z(n2195) );
  ND2SVTX8 U3436 ( .A(n570), .B(n3337), .Z(n1676) );
  ND2SVTX4 U3437 ( .A(n1372), .B(n709), .Z(n2841) );
  EO3SVTX8 U3438 ( .A(n1372), .B(n2176), .C(n3068), .Z(n2842) );
  AO4SVTX6 U3439 ( .A(n2335), .B(n2839), .C(n1083), .D(n2753), .Z(n1372) );
  IVSVTX4 U3440 ( .A(n3571), .Z(n1373) );
  IVSVTX4 U3441 ( .A(n1379), .Z(n1378) );
  ND2SVTX4 U3442 ( .A(n3665), .B(n1821), .Z(n1384) );
  IVSVTX4 U3443 ( .A(n1388), .Z(n2494) );
  IVSVTX12 U3444 ( .A(n1390), .Z(n4138) );
  ND2SVTX8 U3445 ( .A(n2262), .B(n3673), .Z(n1390) );
  AO1CDSVTX6 U3446 ( .A(n1391), .B(n4291), .C(n4189), .D(n4288), .Z(n4270) );
  ND2SVTX4 U3447 ( .A(n1987), .B(n1392), .Z(n1403) );
  IVSVTX12 U3448 ( .A(n1393), .Z(n1419) );
  AO6SVTX8 U3449 ( .A(n2435), .B(n2569), .C(n1418), .Z(n1393) );
  IVSVTX2 U3450 ( .A(n3050), .Z(n1395) );
  AO7ABSVTX4 U3451 ( .A(n3126), .B(n4035), .C(n3391), .Z(n1394) );
  AO6CSVTX6 U3452 ( .A(n3370), .B(n3371), .C(n596), .Z(n1738) );
  ND3SVTX6 U3453 ( .A(n3392), .B(n3391), .C(n482), .Z(n3370) );
  AO7SVTX6 U3454 ( .A(n3788), .B(n3052), .C(n3737), .Z(n3392) );
  ND2SVTX4 U3455 ( .A(n3102), .B(n1395), .Z(n3788) );
  ND2SVTX4 U3456 ( .A(n3056), .B(n3045), .Z(n3390) );
  ND2SVTX4 U3457 ( .A(n2940), .B(n862), .Z(n1399) );
  ND2SVTX4 U3458 ( .A(n1417), .B(n2171), .Z(n1400) );
  IVSVTX4 U3459 ( .A(n3995), .Z(n1401) );
  ND2SVTX4 U3460 ( .A(n524), .B(n3300), .Z(n1402) );
  ND2SVTX8 U3461 ( .A(n1812), .B(n1811), .Z(n1410) );
  IVSVTX4 U3462 ( .A(n2275), .Z(n1413) );
  AO17SVTX8 U3463 ( .A(n1417), .B(n2171), .C(n3995), .D(n1328), .Z(n3299) );
  ND2SVTX8 U3464 ( .A(n2736), .B(n2735), .Z(n1770) );
  IVSVTX4 U3465 ( .A(n1420), .Z(n2407) );
  ND2SVTX6 U3466 ( .A(n1942), .B(n3085), .Z(n3815) );
  AO6SVTX4 U3467 ( .A(n3872), .B(n1426), .C(n1425), .Z(n3822) );
  NR2SVTX4 U3468 ( .A(n928), .B(n3870), .Z(n1426) );
  ND2SVTX4 U3469 ( .A(n3150), .B(n4179), .Z(n3154) );
  AO6SVTX4 U3470 ( .A(n3204), .B(n3201), .C(n3202), .Z(n3155) );
  NR2SVTX8 U3471 ( .A(n1766), .B(n3483), .Z(n1435) );
  EO3SVTX8 U3472 ( .A(n808), .B(n2846), .C(n2168), .Z(n2845) );
  IVSVTX4 U3473 ( .A(n2843), .Z(n1438) );
  ND3ABSVTX8 U3474 ( .A(n1440), .B(n2159), .C(n1439), .Z(n1446) );
  NR2ASVTX6 U3475 ( .A(n4174), .B(n4136), .Z(n1440) );
  AO20SVTX8 U3476 ( .A(n1447), .B(n1446), .C(n4146), .D(n1444), .Z(n4165) );
  IVSVTX4 U3477 ( .A(n4137), .Z(n1447) );
  NR2SVTX4 U3478 ( .A(n3712), .B(n595), .Z(n3709) );
  ENSVTX4 U3479 ( .A(n1450), .B(n2845), .Z(n3484) );
  NR2SVTX4 U3480 ( .A(n2248), .B(n3107), .Z(n1455) );
  NR2SVTX6 U3481 ( .A(n4029), .B(n1464), .Z(n4054) );
  IVSVTX4 U3482 ( .A(n2083), .Z(n1466) );
  EN3SVTX8 U3483 ( .A(n1644), .B(n1939), .C(n1717), .Z(n3460) );
  NR2ASVTX8 U3484 ( .A(n2386), .B(n1475), .Z(n4224) );
  ND2SVTX4 U3485 ( .A(n1476), .B(n1475), .Z(n4225) );
  ND3SVTX8 U3486 ( .A(n3807), .B(n1680), .C(n3806), .Z(n1475) );
  NR2SVTX6 U3487 ( .A(num_i[25]), .B(num_i[29]), .Z(n1477) );
  NR2SVTX6 U3488 ( .A(num_i[26]), .B(num_i[24]), .Z(n1478) );
  AO7ABSVTX4 U3489 ( .A(n1483), .B(n1571), .C(n1578), .Z(n1577) );
  AN3ABCSVTX2 U3490 ( .A(n1482), .B(n3240), .C(n3241), .Z(n3242) );
  B_ND2SVTX2 U3491 ( .A(n3323), .B(n3324), .Z(n4117) );
  NR2ASVTX8 U3492 ( .A(n610), .B(n2964), .Z(n4119) );
  ND2ASVTX8 U3493 ( .A(n604), .B(n3011), .Z(n1488) );
  ND2SVTX6 U3494 ( .A(n1474), .B(n1489), .Z(n1976) );
  ND3SVTX6 U3495 ( .A(n2941), .B(n1292), .C(n1491), .Z(n1492) );
  EO3SVTX8 U3496 ( .A(n2799), .B(n1581), .C(n2934), .Z(n3215) );
  AO7CSVTX8 U3497 ( .A(n1493), .B(n1492), .C(n1490), .Z(n2942) );
  IVSVTX4 U3498 ( .A(n2010), .Z(n2317) );
  B_ND2SVTX2 U3499 ( .A(n3111), .B(n2941), .Z(n1498) );
  IVSVTX4 U3500 ( .A(n1840), .Z(n1839) );
  ND2ASVTX8 U3501 ( .A(n2052), .B(n511), .Z(n1840) );
  ND2SVTX4 U3502 ( .A(n3784), .B(n4009), .Z(n2463) );
  ND3ABSVTX8 U3503 ( .A(n3828), .B(n1870), .C(n1500), .Z(n4009) );
  IVSVTX6 U3504 ( .A(n1502), .Z(n3764) );
  ND3SVTX8 U3505 ( .A(n2358), .B(n3897), .C(n1884), .Z(n3413) );
  NR2SVTX8 U3506 ( .A(n3416), .B(n3415), .Z(n2336) );
  ND3ASVTX6 U3507 ( .A(n2004), .B(n1504), .C(n2003), .Z(n2002) );
  ND2ASVTX8 U3508 ( .A(n1823), .B(n1506), .Z(n1824) );
  ND2SVTX4 U3509 ( .A(n1508), .B(n1512), .Z(n1507) );
  ND2SVTX4 U3510 ( .A(n1816), .B(n1511), .Z(n1509) );
  ND2ASVTX8 U3511 ( .A(n2266), .B(n2180), .Z(n2650) );
  NR2SVTX8 U3512 ( .A(n2329), .B(n2919), .Z(n1516) );
  EO3SVTX8 U3513 ( .A(n1529), .B(n808), .C(n539), .Z(n2917) );
  NR2SVTX4 U3514 ( .A(n579), .B(n2356), .Z(n1519) );
  NR2SVTX2 U3515 ( .A(n1520), .B(n2942), .Z(n2356) );
  NR2SVTX4 U3516 ( .A(n4092), .B(n1554), .Z(n1520) );
  NR2SVTX4 U3517 ( .A(n1644), .B(n1523), .Z(n1522) );
  NR2ASVTX4 U3518 ( .A(n1524), .B(n1525), .Z(n3985) );
  NR2SVTX8 U3519 ( .A(n1740), .B(n1885), .Z(n1525) );
  ND2SVTX8 U3520 ( .A(n1528), .B(n1527), .Z(n1529) );
  ND3SVTX8 U3521 ( .A(n3997), .B(n3996), .C(n1530), .Z(n4025) );
  IVSVTX4 U3522 ( .A(n4066), .Z(n1532) );
  F_IVSVTX1 U3523 ( .A(n2052), .Z(n3846) );
  ND3SVTX8 U3524 ( .A(n548), .B(n2615), .C(n1534), .Z(n2782) );
  EN3SVTX8 U3525 ( .A(n625), .B(n503), .C(n948), .Z(n1906) );
  ND2SVTX6 U3526 ( .A(n2901), .B(n1535), .Z(n3920) );
  ND2SVTX6 U3527 ( .A(n3032), .B(n2865), .Z(n2297) );
  NR2SVTX4 U3528 ( .A(n554), .B(n2364), .Z(n1543) );
  ND2SVTX4 U3529 ( .A(n920), .B(n513), .Z(n1545) );
  AO7CSVTX6 U3530 ( .A(n3311), .B(n3111), .C(n615), .Z(n2875) );
  ND3SVTX6 U3531 ( .A(n1587), .B(n3219), .C(n1548), .Z(n1550) );
  IVSVTX4 U3532 ( .A(n1549), .Z(n1548) );
  ND2ASVTX8 U3533 ( .A(n516), .B(n3215), .Z(n3219) );
  ND2SVTX4 U3534 ( .A(n1553), .B(n1552), .Z(n3457) );
  ND2SVTX4 U3535 ( .A(n4070), .B(n1558), .Z(n1556) );
  IVSVTX4 U3536 ( .A(n1561), .Z(n1558) );
  ND2ASVTX8 U3537 ( .A(n1560), .B(n2827), .Z(n4174) );
  IVSVTX4 U3538 ( .A(n3114), .Z(n1561) );
  ND2SVTX6 U3539 ( .A(n1565), .B(n1563), .Z(n2048) );
  AO7ABSVTX4 U3540 ( .A(n2595), .B(n1022), .C(n2575), .Z(n1563) );
  AO20SVTX8 U3541 ( .A(n1567), .B(n1566), .C(n2245), .D(n2409), .Z(n1565) );
  MUX21NSVTX8 U3542 ( .A(n2517), .B(n635), .S(n1107), .Z(n1566) );
  ND2SVTX4 U3543 ( .A(n1287), .B(n2705), .Z(n1569) );
  IVSVTX4 U3544 ( .A(n4107), .Z(n3057) );
  ND2SVTX8 U3545 ( .A(n1579), .B(n2706), .Z(n2776) );
  ND2SVTX4 U3546 ( .A(n2349), .B(n1715), .Z(n3018) );
  ND2SVTX8 U3547 ( .A(n2557), .B(n2556), .Z(n1580) );
  IVSVTX4 U3548 ( .A(n1580), .Z(n1774) );
  ND2SVTX8 U3549 ( .A(n2793), .B(n2792), .Z(n2934) );
  ND2SVTX4 U3550 ( .A(n3165), .B(n2869), .Z(n2929) );
  EO3SVTX8 U3551 ( .A(n622), .B(n2790), .C(n2791), .Z(n2937) );
  ND3SVTX2 U3552 ( .A(n2399), .B(n485), .C(n1690), .Z(n3884) );
  BFSVTX10 U3553 ( .A(n1090), .Z(n2240) );
  IVSVTX12 U3554 ( .A(n2246), .Z(n2582) );
  ND3ABSVTX6 U3555 ( .A(num_i[24]), .B(num_i[25]), .C(n2479), .Z(n2482) );
  IVSVTX4 U3556 ( .A(n3824), .Z(n3819) );
  NR2ASVTX6 U3557 ( .A(n1268), .B(n519), .Z(n1598) );
  EN3SVTX8 U3558 ( .A(n2888), .B(n508), .C(n626), .Z(n2316) );
  IVSVTX4 U3559 ( .A(n4159), .Z(n3132) );
  AO7SVTX4 U3560 ( .A(n502), .B(n627), .C(n1741), .Z(n2404) );
  NR3ABSVTX8 U3561 ( .A(n2664), .B(n1598), .C(n2342), .Z(n2725) );
  OR2SVTX4 U3562 ( .A(n550), .B(n2561), .Z(n2504) );
  NR2SVTX6 U3563 ( .A(n3928), .B(n3802), .Z(n3803) );
  NR2SVTX2 U3564 ( .A(n4073), .B(n506), .Z(n4131) );
  EOSVTX8 U3565 ( .A(n1025), .B(n684), .Z(n2068) );
  AO7SVTX4 U3566 ( .A(n3185), .B(n4037), .C(n3176), .Z(n3177) );
  ND2SVTX2 U3567 ( .A(n2760), .B(n1268), .Z(n2758) );
  IVSVTX12 U3568 ( .A(n2561), .Z(n1756) );
  NR2SVTX4 U3569 ( .A(n2526), .B(n2525), .Z(n2530) );
  ND3SVTX8 U3570 ( .A(n3583), .B(n3626), .C(n1980), .Z(n2976) );
  IVSVTX4 U3571 ( .A(n1748), .Z(n1882) );
  EN3SVTX8 U3572 ( .A(n1025), .B(n1967), .C(n2971), .Z(n2138) );
  ENSVTX8 U3573 ( .A(n1939), .B(n1940), .Z(n3503) );
  AN2SVTX4 U3574 ( .A(n2812), .B(n1419), .Z(n2710) );
  ND2ASVTX8 U3575 ( .A(n2542), .B(n2541), .Z(n2110) );
  NR2ASVTX6 U3576 ( .A(n3510), .B(n3509), .Z(n3511) );
  EN3SVTX8 U3577 ( .A(n643), .B(n1042), .C(n1973), .Z(n1979) );
  AO2SVTX8 U3578 ( .A(n2786), .B(n2777), .C(n506), .D(n1679), .Z(n2417) );
  ND2SVTX6 U3579 ( .A(n3343), .B(n3344), .Z(n3387) );
  IVSVTX12 U3580 ( .A(n1607), .Z(n2587) );
  ND2ASVTX8 U3581 ( .A(n1107), .B(n1297), .Z(n1607) );
  NR2SVTX4 U3582 ( .A(n1611), .B(n3686), .Z(n3547) );
  IVSVTX10 U3583 ( .A(n2172), .Z(n2171) );
  IVSVTX4 U3584 ( .A(n1613), .Z(n2403) );
  ND2SVTX4 U3585 ( .A(n1022), .B(n1872), .Z(n1613) );
  AO4SVTX8 U3586 ( .A(n2838), .B(n2839), .C(n1083), .D(n2632), .Z(n2888) );
  ND2SVTX4 U3587 ( .A(n3508), .B(n3519), .Z(n1615) );
  AO1CDSVTX8 U3588 ( .A(n1896), .B(n2234), .C(n1596), .D(n3409), .Z(n1841) );
  AO3SVTX6 U3589 ( .A(n1698), .B(n4023), .C(n2446), .D(n1636), .Z(n3651) );
  EN3SVTX8 U3590 ( .A(n2945), .B(n1571), .C(n1728), .Z(n2951) );
  ND2SVTX4 U3591 ( .A(n4015), .B(n1616), .Z(n4016) );
  ND2SVTX4 U3592 ( .A(n4014), .B(n4013), .Z(n1616) );
  ND3SVTX8 U3593 ( .A(n3991), .B(n2441), .C(n3992), .Z(n1670) );
  AN3SVTX6 U3594 ( .A(n514), .B(n575), .C(n4021), .Z(n2430) );
  AO7ABSVTX4 U3595 ( .A(n686), .B(n684), .C(n1620), .Z(n3504) );
  ND2SVTX4 U3596 ( .A(n1621), .B(n1042), .Z(n1620) );
  NR2SVTX4 U3597 ( .A(n684), .B(n686), .Z(n1622) );
  EO3SVTX8 U3598 ( .A(n659), .B(n686), .C(n1042), .Z(n3075) );
  NR2SVTX8 U3599 ( .A(n2712), .B(n2711), .Z(n2713) );
  NR2ASVTX2 U3600 ( .A(n2579), .B(n2503), .Z(n2580) );
  NR2SVTX4 U3601 ( .A(n3311), .B(n2378), .Z(n3161) );
  NR2SVTX4 U3602 ( .A(n2391), .B(n2282), .Z(n2390) );
  AO7SVTX6 U3603 ( .A(n2740), .B(n2739), .C(n2738), .Z(n2741) );
  AO7SVTX4 U3604 ( .A(n1704), .B(n1703), .C(n2217), .Z(n4067) );
  AO7SVTX4 U3605 ( .A(n428), .B(n1481), .C(n1939), .Z(n1813) );
  AO7SVTX6 U3606 ( .A(n3728), .B(n1740), .C(n4066), .Z(n3729) );
  NR2SVTX4 U3607 ( .A(n4274), .B(n1678), .Z(n4088) );
  ND4ABSVTX8 U3608 ( .A(n3894), .B(n524), .C(n3901), .D(n3900), .Z(n3902) );
  ND2SVTX4 U3609 ( .A(n530), .B(n3481), .Z(n3482) );
  IVSVTX4 U3610 ( .A(n1630), .Z(n3947) );
  AO7ABSVTX4 U3611 ( .A(n441), .B(n814), .C(n3848), .Z(n1754) );
  ND2SVTX4 U3612 ( .A(n626), .B(n1631), .Z(n2146) );
  IVSVTX4 U3613 ( .A(n1938), .Z(n1631) );
  NR2SVTX4 U3614 ( .A(n3079), .B(n1647), .Z(n1938) );
  ND2SVTX2 U3615 ( .A(n1661), .B(n3474), .Z(n3475) );
  ND3ASVTX4 U3616 ( .A(n516), .B(n3310), .C(n1719), .Z(n3246) );
  ND2SVTX4 U3617 ( .A(n2606), .B(n2607), .Z(n2700) );
  EN3SVTX6 U3618 ( .A(n616), .B(n1764), .C(n1789), .Z(n3053) );
  AO7SVTX6 U3619 ( .A(n2935), .B(n2934), .C(n2933), .Z(n2011) );
  AO4SVTX8 U3620 ( .A(n918), .B(n1721), .C(n2902), .D(n632), .Z(n2993) );
  B_ND2SVTX2 U3621 ( .A(n2424), .B(n3658), .Z(n2439) );
  ND2SVTX4 U3622 ( .A(n514), .B(n3019), .Z(n2828) );
  MUX21NSVTX4 U3623 ( .A(n3530), .B(n373), .S(n3484), .Z(n2063) );
  IVSVTX12 U3624 ( .A(n836), .Z(n2971) );
  AO7NSVTX4 U3625 ( .A(n3766), .B(n3885), .C(n3853), .Z(n2405) );
  ND2SVTX4 U3626 ( .A(n3613), .B(n3180), .Z(n3183) );
  IVSVTX4 U3627 ( .A(n3616), .Z(n1639) );
  AO7ABSVTX4 U3628 ( .A(n3067), .B(n3068), .C(n3069), .Z(n3459) );
  ND4SVTX4 U3629 ( .A(n3808), .B(n3820), .C(n924), .D(n3930), .Z(n1640) );
  IVSVTX4 U3630 ( .A(n2014), .Z(n1643) );
  AO7ABSVTX8 U3631 ( .A(n2779), .B(n3111), .C(n2778), .Z(n2780) );
  ND4ABCSVTX8 U3632 ( .A(n1858), .B(n2572), .C(n2126), .D(n2245), .Z(n2697) );
  NR2SVTX4 U3633 ( .A(n1649), .B(n2757), .Z(n2116) );
  ND2ASVTX8 U3634 ( .A(n3065), .B(n1826), .Z(n3066) );
  NR2SVTX4 U3635 ( .A(n2636), .B(n2613), .Z(n2686) );
  ND2SVTX4 U3636 ( .A(n633), .B(n2705), .Z(n2706) );
  NR2SVTX4 U3637 ( .A(n4208), .B(n4205), .Z(n4210) );
  AN2SVTX4 U3638 ( .A(n3632), .B(n3631), .Z(n2458) );
  IVSVTX12 U3639 ( .A(n4138), .Z(n2351) );
  NR4SVTX8 U3640 ( .A(n2743), .B(n2728), .C(n2088), .D(n2087), .Z(n2263) );
  ND2ASVTX8 U3641 ( .A(n1807), .B(n2995), .Z(n3544) );
  ND3ABSVTX8 U3642 ( .A(n1473), .B(n1871), .C(n1852), .Z(n4023) );
  AO7ABSVTX8 U3643 ( .A(n2238), .B(n1872), .C(n1916), .Z(n2334) );
  ND2SVTX6 U3644 ( .A(n1360), .B(n2676), .Z(n2663) );
  IVSVTX4 U3645 ( .A(n3861), .Z(n3862) );
  ND2ASVTX8 U3646 ( .A(n844), .B(n2197), .Z(n3736) );
  ND2ASVTX8 U3647 ( .A(n2306), .B(n2048), .Z(n2305) );
  NR2SVTX2 U3648 ( .A(n2370), .B(n2784), .Z(n2785) );
  AO8SVTX6 U3649 ( .A(n3438), .B(n3445), .C(n3444), .D(n2259), .Z(n2436) );
  EO3SVTX6 U3650 ( .A(n625), .B(n1339), .C(n3311), .Z(n3096) );
  ENSVTX8 U3651 ( .A(n479), .B(n2140), .Z(n1694) );
  AO17SVTX4 U3652 ( .A(n622), .B(n3145), .C(n3144), .D(n1667), .Z(n2212) );
  ND2SVTX4 U3653 ( .A(n2456), .B(n3012), .Z(n4175) );
  IVSVTX4 U3654 ( .A(n4225), .Z(n1668) );
  ND2ASVTX8 U3655 ( .A(n3688), .B(n3560), .Z(n4258) );
  F_ND3SVTX2 U3656 ( .A(n594), .B(n392), .C(n578), .Z(n2004) );
  AO7ABSVTX8 U3657 ( .A(n2624), .B(n1768), .C(n1672), .Z(n2661) );
  ND3SVTX8 U3658 ( .A(n4028), .B(n4027), .C(n4026), .Z(n1673) );
  ND2SVTX6 U3659 ( .A(n4295), .B(n1933), .Z(n3910) );
  ND3SVTX8 U3660 ( .A(n1857), .B(n2561), .C(n2551), .Z(n1904) );
  ND2ASVTX8 U3661 ( .A(n2127), .B(n2487), .Z(n2551) );
  AO7SVTX8 U3662 ( .A(n1914), .B(n4216), .C(n4213), .Z(n4297) );
  IVSVTX4 U3663 ( .A(n2961), .Z(n2959) );
  EO3SVTX8 U3664 ( .A(n686), .B(n911), .C(n1618), .Z(n2890) );
  BFSVTX6 U3665 ( .A(n4268), .Z(n1678) );
  EO3SVTX8 U3666 ( .A(n506), .B(n1855), .C(n2786), .Z(n2010) );
  AO1ABSVTX8 U3667 ( .A(n697), .B(n2109), .C(n2106), .D(n2104), .Z(n1680) );
  ND2SVTX4 U3668 ( .A(n1681), .B(n3041), .Z(n3054) );
  AO17SVTX8 U3669 ( .A(n2607), .B(n2606), .C(n2612), .D(n2605), .Z(n2608) );
  IVSVTX4 U3670 ( .A(n1682), .Z(n2406) );
  AO3SVTX8 U3671 ( .A(n4214), .B(n3910), .C(n3909), .D(n2434), .Z(n4221) );
  MUX21NSVTX2 U3672 ( .A(n3837), .B(n3836), .S(n4014), .Z(n3838) );
  IVSVTX2 U3673 ( .A(n3746), .Z(n3747) );
  AO6SVTX4 U3674 ( .A(n3755), .B(n3756), .C(n495), .Z(n1683) );
  ND2SVTX4 U3675 ( .A(n2149), .B(n623), .Z(n3887) );
  ND2SVTX4 U3676 ( .A(n2478), .B(n2518), .Z(n2479) );
  NR2SVTX4 U3677 ( .A(n3135), .B(n526), .Z(n3131) );
  NR2SVTX4 U3678 ( .A(n3124), .B(n3123), .Z(n3135) );
  ND3ASVTX8 U3679 ( .A(n3698), .B(n1749), .C(n1832), .Z(n1817) );
  NR2SVTX4 U3680 ( .A(n2599), .B(n650), .Z(n1687) );
  BFSVTX1 U3681 ( .A(n4257), .Z(n1688) );
  IVSVTX2 U3682 ( .A(n2374), .Z(n3882) );
  AO7ABSVTX4 U3683 ( .A(n1689), .B(n974), .C(n3881), .Z(n3883) );
  ND2SVTX4 U3684 ( .A(n1692), .B(n1691), .Z(n1799) );
  IVSVTX4 U3685 ( .A(n1693), .Z(n3335) );
  ND2SVTX6 U3686 ( .A(n3591), .B(n3590), .Z(n3584) );
  ND3SVTX6 U3687 ( .A(n3337), .B(n1705), .C(n570), .Z(n3319) );
  IVSVTX4 U3688 ( .A(n3780), .Z(n1696) );
  NR2ASVTX6 U3689 ( .A(n3311), .B(n1700), .Z(n2054) );
  NR3SVTX8 U3690 ( .A(n3283), .B(n1634), .C(n2731), .Z(n2732) );
  EN3SVTX8 U3691 ( .A(n1764), .B(n623), .C(n3272), .Z(n3102) );
  EOSVTX4 U3692 ( .A(n4228), .B(n4227), .Z(rslt_o[11]) );
  CTIVSVTX4 U3693 ( .A(n2168), .Z(n1710) );
  AO7SVTX2 U3694 ( .A(n4298), .B(n1720), .C(n1757), .Z(n4299) );
  BFSVTX6 U3695 ( .A(n3815), .Z(n3930) );
  ND3SVTX8 U3696 ( .A(n2756), .B(n2253), .C(n2116), .Z(n2117) );
  IVSVTX8 U3697 ( .A(n2111), .Z(n1871) );
  NR3ABSVTX8 U3698 ( .A(n2528), .B(n2509), .C(n2366), .Z(n2487) );
  IVSVTX8 U3699 ( .A(n1712), .Z(n2111) );
  NR3ASVTX6 U3700 ( .A(n553), .B(n2527), .C(n2033), .Z(n2529) );
  NR3ASVTX6 U3701 ( .A(n3402), .B(n3399), .C(n3407), .Z(n1846) );
  ND3SVTX6 U3702 ( .A(n2379), .B(n2018), .C(n2981), .Z(n2381) );
  NR2SVTX4 U3703 ( .A(n554), .B(n1768), .Z(n1708) );
  ND2ASVTX8 U3704 ( .A(n1711), .B(n2976), .Z(n3960) );
  AO4SVTX8 U3705 ( .A(n2864), .B(n2863), .C(n3566), .D(n2372), .Z(n1712) );
  NR2SVTX4 U3706 ( .A(n3182), .B(n1713), .Z(n3199) );
  NR2SVTX2 U3707 ( .A(n1892), .B(n3272), .Z(n2968) );
  IVSVTX4 U3708 ( .A(n3053), .Z(n1714) );
  BFSVTX6 U3709 ( .A(n1268), .Z(n1717) );
  AO7SVTX6 U3710 ( .A(n3932), .B(n3931), .C(n3929), .Z(n1718) );
  BFSVTX1 U3711 ( .A(n4224), .Z(n1720) );
  BFSVTX1 U3712 ( .A(n4260), .Z(n1722) );
  IVSVTX4 U3713 ( .A(n2316), .Z(n3449) );
  ND2ASVTX8 U3714 ( .A(n2222), .B(n3299), .Z(n4167) );
  ND2SVTX4 U3715 ( .A(n1726), .B(n1725), .Z(n4123) );
  ND2SVTX4 U3716 ( .A(n2978), .B(n2130), .Z(n1921) );
  ND2SVTX4 U3717 ( .A(n1733), .B(n3269), .Z(n2214) );
  IVSVTX2 U3718 ( .A(n4270), .Z(n1736) );
  NR2SVTX2 U3719 ( .A(n4273), .B(n4272), .Z(n1737) );
  IVSVTX6 U3720 ( .A(n1090), .Z(n1937) );
  NR2ASVTX6 U3721 ( .A(n3365), .B(n1738), .Z(n3313) );
  IVSVTX8 U3722 ( .A(n2864), .Z(n2016) );
  ND3SVTX8 U3723 ( .A(n1336), .B(n521), .C(n2661), .Z(n2655) );
  NR4ABSVTX8 U3724 ( .A(n1343), .B(n2247), .C(n3470), .D(n3905), .Z(n2249) );
  EN3SVTX8 U3725 ( .A(n3065), .B(n1939), .C(n612), .Z(n3551) );
  NR2ASVTX6 U3726 ( .A(n644), .B(n586), .Z(n3851) );
  AO6CSVTX4 U3727 ( .A(n2225), .B(n4201), .C(n4200), .Z(n4198) );
  BFSVTX6 U3728 ( .A(n2489), .Z(n1744) );
  NR2SVTX4 U3729 ( .A(n3190), .B(n3189), .Z(n3192) );
  ND3ABSVTX8 U3730 ( .A(n1022), .B(n1360), .C(n2654), .Z(n2656) );
  IVSVTX2 U3731 ( .A(n2804), .Z(n2802) );
  ENSVTX8 U3732 ( .A(n4206), .B(n1802), .Z(rslt_o[24]) );
  ND2SVTX4 U3733 ( .A(n2065), .B(n1747), .Z(n2062) );
  ND2SVTX4 U3734 ( .A(n543), .B(n1777), .Z(n2251) );
  NR2SVTX4 U3735 ( .A(n1818), .B(n1833), .Z(n1749) );
  AO7ABSVTX8 U3736 ( .A(n2199), .B(n2820), .C(n1798), .Z(n1801) );
  AN2SVTX4 U3737 ( .A(n1903), .B(n637), .Z(n2607) );
  AO5SVTX6 U3738 ( .A(n615), .B(n2387), .C(n2954), .Z(n2950) );
  IVSVTX4 U3739 ( .A(n2950), .Z(n2953) );
  BFSVTX6 U3740 ( .A(num_i[14]), .Z(n1755) );
  AO6SVTX6 U3741 ( .A(n2482), .B(n2481), .C(n2480), .Z(n2485) );
  BFSVTX1 U3742 ( .A(n4225), .Z(n1757) );
  ND2ASVTX8 U3743 ( .A(n3001), .B(n1758), .Z(n3590) );
  NR2ASVTX6 U3744 ( .A(n2657), .B(n1761), .Z(n1957) );
  ND2SVTX6 U3745 ( .A(n2423), .B(n3965), .Z(n3326) );
  IVSVTX4 U3746 ( .A(n3326), .Z(n1787) );
  F_EOSVTX2 U3747 ( .A(n2784), .B(n541), .Z(n1788) );
  ND2SVTX4 U3748 ( .A(n1793), .B(n1792), .Z(n3007) );
  EN3SVTX8 U3749 ( .A(n3283), .B(n1397), .C(n2151), .Z(n1794) );
  ND2SVTX4 U3750 ( .A(n4047), .B(n1795), .Z(n4049) );
  ND2ASVTX8 U3751 ( .A(n3653), .B(n2111), .Z(n1796) );
  ND2SVTX8 U3752 ( .A(n2862), .B(n2861), .Z(n3653) );
  NR2ASVTX6 U3753 ( .A(n1107), .B(n1323), .Z(n1797) );
  ND2SVTX4 U3754 ( .A(n1656), .B(n2048), .Z(n2615) );
  AO7SVTX6 U3755 ( .A(n1800), .B(n1801), .C(n1799), .Z(n2179) );
  AO7SVTX8 U3756 ( .A(n4273), .B(n4272), .C(n4270), .Z(n2225) );
  AO6SVTX8 U3757 ( .A(n4221), .B(n4054), .C(n4053), .Z(n4272) );
  AO6SVTX4 U3758 ( .A(n2225), .B(n1804), .C(n1803), .Z(n1802) );
  NR2SVTX4 U3759 ( .A(n4166), .B(n4205), .Z(n1804) );
  IVSVTX4 U3760 ( .A(n2753), .Z(n2632) );
  ND2SVTX4 U3761 ( .A(n603), .B(n2996), .Z(n3539) );
  AO7SVTX8 U3762 ( .A(n3544), .B(n1699), .C(n3539), .Z(n3586) );
  ND2SVTX8 U3763 ( .A(n3594), .B(n2402), .Z(n3965) );
  ND2SVTX4 U3764 ( .A(n428), .B(n1481), .Z(n1814) );
  AO21DSVTX8 U3765 ( .A(n1819), .B(n3650), .C(n1817), .D(n522), .Z(n2102) );
  NR2SVTX4 U3766 ( .A(n524), .B(n3700), .Z(n1819) );
  AO7SVTX6 U3767 ( .A(n3716), .B(n2413), .C(n566), .Z(n4230) );
  NR3ABSVTX8 U3768 ( .A(n4066), .B(n3715), .C(n1820), .Z(n2413) );
  IVSVTX4 U3769 ( .A(n2115), .Z(n2628) );
  ND2SVTX8 U3770 ( .A(n486), .B(n3742), .Z(n4159) );
  ND2SVTX8 U3771 ( .A(n3789), .B(n3172), .Z(n3742) );
  ND2SVTX4 U3772 ( .A(n1827), .B(n2240), .Z(n3063) );
  IVSVTX4 U3773 ( .A(n1829), .Z(n3964) );
  ND2SVTX4 U3774 ( .A(n2443), .B(n2396), .Z(n3966) );
  NR2SVTX4 U3775 ( .A(n1830), .B(n1829), .Z(n2396) );
  ND3SVTX6 U3776 ( .A(n2190), .B(n491), .C(n3722), .Z(n1829) );
  ND2SVTX4 U3777 ( .A(n3965), .B(n744), .Z(n2443) );
  IVSVTX4 U3778 ( .A(n3650), .Z(n1831) );
  AO7SVTX4 U3779 ( .A(n1972), .B(n2129), .C(n728), .Z(n1836) );
  ND2SVTX4 U3780 ( .A(n1937), .B(n543), .Z(n3672) );
  AO7CSVTX6 U3781 ( .A(n1850), .B(n1740), .C(n3417), .Z(n1901) );
  ND2SVTX8 U3782 ( .A(n1796), .B(n528), .Z(n2014) );
  IVSVTX4 U3783 ( .A(n2787), .Z(n1855) );
  ND2SVTX6 U3784 ( .A(n2490), .B(n2406), .Z(n1857) );
  IVSVTX4 U3785 ( .A(n1857), .Z(n1858) );
  ND2SVTX6 U3786 ( .A(n1857), .B(n2561), .Z(n2552) );
  NR2SVTX4 U3787 ( .A(n3261), .B(n2135), .Z(n3262) );
  ND3ASVTX6 U3788 ( .A(n3297), .B(n977), .C(n2361), .Z(n3300) );
  ND2ASVTX8 U3789 ( .A(n918), .B(n1859), .Z(n2783) );
  ND2SVTX8 U3790 ( .A(n2782), .B(n2783), .Z(n3032) );
  ND2SVTX4 U3791 ( .A(n1866), .B(n2117), .Z(n1873) );
  ND3SVTX8 U3792 ( .A(n2725), .B(n2724), .C(n2713), .Z(n1945) );
  ND2SVTX4 U3793 ( .A(n2577), .B(n2486), .Z(n2480) );
  ND2SVTX4 U3794 ( .A(n2814), .B(n1686), .Z(n3827) );
  ND3SVTX8 U3795 ( .A(n1872), .B(n2636), .C(n2355), .Z(n2649) );
  ND2SVTX8 U3796 ( .A(n1886), .B(n1887), .Z(n3280) );
  NR2SVTX8 U3797 ( .A(n1890), .B(n4224), .Z(n1933) );
  IVSVTX4 U3798 ( .A(n1890), .Z(n4294) );
  IVSVTX4 U3799 ( .A(n4293), .Z(n1891) );
  ND2SVTX4 U3800 ( .A(n2329), .B(n2919), .Z(n3763) );
  ND3SVTX8 U3801 ( .A(n1287), .B(n1895), .C(n2560), .Z(n2811) );
  IVSVTX4 U3802 ( .A(n4171), .Z(n3383) );
  IVSVTX4 U3803 ( .A(n1902), .Z(n4000) );
  IVSVTX4 U3804 ( .A(n1907), .Z(n2901) );
  EN3SVTX8 U3805 ( .A(n544), .B(n547), .C(n3078), .Z(n2168) );
  ND2SVTX4 U3806 ( .A(n533), .B(n1909), .Z(n3402) );
  ND2SVTX4 U3807 ( .A(n4030), .B(n415), .Z(n3398) );
  ND3SVTX6 U3808 ( .A(n2528), .B(n1913), .C(n460), .Z(n2547) );
  IVSVTX12 U3809 ( .A(n2657), .Z(n2678) );
  AO6SVTX8 U3810 ( .A(n2204), .B(n2205), .C(n2203), .Z(n3789) );
  IVSVTX4 U3811 ( .A(n3171), .Z(n3792) );
  EN3SVTX8 U3812 ( .A(n2375), .B(n1851), .C(n1791), .Z(n3957) );
  ND2ASVTX8 U3813 ( .A(n1923), .B(n3027), .Z(n3245) );
  F_ENSVTX2 U3814 ( .A(n1924), .B(n2392), .Z(n3121) );
  F_EOSVTX2 U3815 ( .A(n2789), .B(n2720), .Z(n1924) );
  ND2SVTX6 U3816 ( .A(n1933), .B(n4297), .Z(n3909) );
  NR2SVTX4 U3817 ( .A(n3779), .B(n3866), .Z(n3782) );
  NR2SVTX4 U3818 ( .A(n1935), .B(n3781), .Z(n2076) );
  NR2SVTX4 U3819 ( .A(n2019), .B(n584), .Z(n3781) );
  IVSVTX8 U3820 ( .A(num_i[24]), .Z(n2133) );
  ENSVTX8 U3821 ( .A(n1090), .B(n3079), .Z(n1940) );
  AO7SVTX4 U3822 ( .A(n1938), .B(n964), .C(n2147), .Z(n3082) );
  AO7SVTX6 U3823 ( .A(n2744), .B(n1945), .C(n1984), .Z(n2262) );
  ND2SVTX1 U3824 ( .A(n1946), .B(n2102), .Z(n4240) );
  ND2ASVTX8 U3825 ( .A(n2905), .B(n2198), .Z(n2360) );
  IVSVTX4 U3826 ( .A(n1947), .Z(n1948) );
  ND2SVTX8 U3827 ( .A(n1954), .B(n1955), .Z(n4018) );
  ND2SVTX4 U3828 ( .A(n3287), .B(n3433), .Z(n1959) );
  IVSVTX4 U3829 ( .A(n3981), .Z(n3984) );
  ND2SVTX8 U3830 ( .A(n4022), .B(n3845), .Z(n3948) );
  ND2SVTX8 U3831 ( .A(n2860), .B(n2859), .Z(n3845) );
  ND2SVTX2 U3832 ( .A(n1975), .B(n2854), .Z(n2853) );
  ND2SVTX8 U3833 ( .A(n2346), .B(n3948), .Z(n2234) );
  NR2SVTX8 U3834 ( .A(n1766), .B(n3483), .Z(n3531) );
  IVSVTX4 U3835 ( .A(n4271), .Z(n4197) );
  ND2SVTX6 U3836 ( .A(n3266), .B(n3265), .Z(n3002) );
  AO6SVTX4 U3837 ( .A(n3303), .B(n3304), .C(n3308), .Z(n1988) );
  NR2SVTX4 U3838 ( .A(n2248), .B(n3314), .Z(n1989) );
  NR2SVTX4 U3839 ( .A(n4007), .B(n4004), .Z(n1991) );
  NR2ASVTX6 U3840 ( .A(n1993), .B(n1992), .Z(n4010) );
  IVSVTX4 U3841 ( .A(n2416), .Z(n1992) );
  ND2SVTX8 U3842 ( .A(n3640), .B(n3641), .Z(n4014) );
  ND2ASVTX6 U3843 ( .A(n3289), .B(n3889), .Z(n3745) );
  ND2SVTX6 U3844 ( .A(n1996), .B(n2677), .Z(n1995) );
  IVSVTX4 U3845 ( .A(n3413), .Z(n1998) );
  NR2SVTX4 U3846 ( .A(n2077), .B(n587), .Z(n2001) );
  IVSVTX4 U3847 ( .A(n4144), .Z(n2003) );
  ND2SVTX8 U3848 ( .A(n2196), .B(n2006), .Z(n3619) );
  ND2SVTX6 U3849 ( .A(n2066), .B(n2008), .Z(n2007) );
  ND2SVTX8 U3850 ( .A(n2011), .B(n2010), .Z(n4068) );
  BFSVTX6 U3851 ( .A(n4068), .Z(n2009) );
  AO7SVTX4 U3852 ( .A(n3068), .B(n3067), .C(n687), .Z(n3069) );
  IVSVTX12 U3853 ( .A(n542), .Z(n3311) );
  NR2ASVTX2 U3854 ( .A(n2930), .B(n3035), .Z(n4140) );
  IVSVTX2 U3855 ( .A(n3576), .Z(n3577) );
  AO7SVTX6 U3856 ( .A(n2017), .B(n537), .C(n3068), .Z(n3058) );
  EN3SVTX8 U3857 ( .A(n808), .B(n502), .C(n3068), .Z(n3089) );
  AO6SVTX4 U3858 ( .A(n2025), .B(n2024), .C(n3336), .Z(n2023) );
  NR2SVTX4 U3859 ( .A(n3976), .B(n3975), .Z(n3978) );
  ND2SVTX4 U3860 ( .A(n2760), .B(n2032), .Z(n2264) );
  IVSVTX4 U3861 ( .A(n659), .Z(n2032) );
  ND2SVTX6 U3862 ( .A(n2313), .B(n2486), .Z(n2526) );
  NR2SVTX6 U3863 ( .A(num_i[18]), .B(num_i[16]), .Z(n2313) );
  ND3ABSVTX8 U3864 ( .A(num_i[19]), .B(num_i[30]), .C(n639), .Z(n2033) );
  ND2SVTX4 U3865 ( .A(n3067), .B(n684), .Z(n3287) );
  NR2SVTX4 U3866 ( .A(n3675), .B(n3678), .Z(n2034) );
  NR2ASVTX6 U3867 ( .A(n2035), .B(n3534), .Z(n3678) );
  NR2SVTX8 U3868 ( .A(n2043), .B(n2039), .Z(n2038) );
  ND4ABSVTX6 U3869 ( .A(n3258), .B(n4073), .C(n2046), .D(n2045), .Z(n2044) );
  ND3SVTX4 U3870 ( .A(n3257), .B(n2135), .C(n2345), .Z(n2045) );
  AO1CDSVTX6 U3871 ( .A(n3257), .B(n4167), .C(n2174), .D(n2173), .Z(n2046) );
  ND2SVTX4 U3872 ( .A(n1494), .B(n466), .Z(n2053) );
  ND2SVTX4 U3873 ( .A(n2009), .B(n3219), .Z(n2056) );
  ND2SVTX4 U3874 ( .A(n548), .B(n2143), .Z(n2319) );
  ND2SVTX4 U3875 ( .A(n3114), .B(n3115), .Z(n3119) );
  NR2ASVTX6 U3876 ( .A(n2941), .B(n2797), .Z(n2058) );
  NR2ASVTX8 U3877 ( .A(n543), .B(n2069), .Z(n3440) );
  AO6CSVTX8 U3878 ( .A(n2750), .B(n1150), .C(n2749), .Z(n3441) );
  ND2ASVTX8 U3879 ( .A(n543), .B(n2069), .Z(n3439) );
  IVSVTX4 U3880 ( .A(n2107), .Z(n2073) );
  ND2SVTX4 U3881 ( .A(n3781), .B(n2075), .Z(n2074) );
  ND2SVTX4 U3882 ( .A(n3629), .B(n3628), .Z(n3780) );
  NR2SVTX8 U3883 ( .A(n2909), .B(n2908), .Z(n2077) );
  IVSVTX4 U3884 ( .A(n2351), .Z(n3854) );
  AO1ABSVTX6 U3885 ( .A(n2351), .B(n2080), .C(n3892), .D(n2079), .Z(n2229) );
  IVSVTX4 U3886 ( .A(n2907), .Z(n2089) );
  NR2ASVTX6 U3887 ( .A(n2092), .B(n2017), .Z(n4004) );
  ND2SVTX4 U3888 ( .A(n2810), .B(n2811), .Z(n2375) );
  AO20SVTX8 U3889 ( .A(n2097), .B(n2094), .C(n3268), .D(n1660), .Z(n2093) );
  ND2SVTX4 U3890 ( .A(n3782), .B(n2374), .Z(n2108) );
  ND2SVTX4 U3891 ( .A(n485), .B(n3782), .Z(n2107) );
  ND2SVTX8 U3892 ( .A(n3719), .B(n3795), .Z(n3928) );
  IVSVTX4 U3893 ( .A(n2117), .Z(n2767) );
  AO6SVTX4 U3894 ( .A(n640), .B(num_i[25]), .C(num_i[27]), .Z(n2522) );
  ENSVTX4 U3895 ( .A(n2225), .B(n4202), .Z(rslt_o[19]) );
  NR4ABCSVTX6 U3896 ( .A(n3221), .B(n3948), .C(n3219), .D(n3214), .Z(n2124) );
  ND2SVTX8 U3897 ( .A(n2540), .B(n2620), .Z(n2570) );
  EN3SVTX8 U3898 ( .A(n1644), .B(n620), .C(n503), .Z(n3958) );
  ND2ASVTX8 U3899 ( .A(n3566), .B(n2131), .Z(n3656) );
  IVSVTX4 U3900 ( .A(n2372), .Z(n2131) );
  AO5SVTX8 U3901 ( .A(n627), .B(n2137), .C(n2848), .Z(n2854) );
  NR2SVTX4 U3902 ( .A(n1030), .B(n2971), .Z(n2141) );
  NR2ASVTX6 U3903 ( .A(n1882), .B(n3283), .Z(n2148) );
  ND2ASVTX6 U3904 ( .A(n579), .B(n558), .Z(n2161) );
  ND2SVTX6 U3905 ( .A(n2939), .B(n2317), .Z(n2936) );
  ND2SVTX4 U3906 ( .A(n2841), .B(n2840), .Z(n2846) );
  AO8ASVTX6 U3907 ( .A(n3233), .B(n3243), .C(n2090), .D(n3242), .Z(n2175) );
  IVSVTX4 U3908 ( .A(n2179), .Z(n2178) );
  IVSVTX6 U3909 ( .A(n513), .Z(n2294) );
  ND4SVTX4 U3910 ( .A(n4094), .B(n2345), .C(n4091), .D(n2181), .Z(n4095) );
  NR2SVTX6 U3911 ( .A(num_i[9]), .B(num_i[8]), .Z(n2472) );
  AO8DSVTX6 U3912 ( .A(n2206), .B(n1658), .C(n3983), .D(n4138), .Z(n2429) );
  EN3SVTX8 U3913 ( .A(n3122), .B(n2781), .C(n2778), .Z(n3212) );
  ND3ABSVTX8 U3914 ( .A(n2219), .B(n2218), .C(n433), .Z(n2217) );
  NR2SVTX8 U3915 ( .A(num_i[22]), .B(num_i[23]), .Z(n2220) );
  AO6CSVTX8 U3916 ( .A(n2225), .B(n4194), .C(n4207), .Z(n4187) );
  AO6SVTX4 U3917 ( .A(n2225), .B(n4088), .C(n4087), .Z(n4089) );
  AO4SVTX6 U3918 ( .A(n2629), .B(n2364), .C(n555), .D(n2294), .Z(n2238) );
  ND2ASVTX8 U3919 ( .A(n3088), .B(n3061), .Z(n3817) );
  BFSVTX6 U3920 ( .A(n2582), .Z(n2245) );
  ND2ASVTX8 U3921 ( .A(n546), .B(n2200), .Z(n3796) );
  IVSVTX4 U3922 ( .A(n2254), .Z(n2253) );
  ND2ASVTX8 U3923 ( .A(n2991), .B(n2283), .Z(n3588) );
  AO7SVTX6 U3924 ( .A(n622), .B(n2791), .C(n2790), .Z(n2792) );
  EO3SVTX8 U3925 ( .A(n2255), .B(n944), .C(n2788), .Z(n2791) );
  NR2SVTX8 U3926 ( .A(n895), .B(n2257), .Z(n2652) );
  ND2ASVTX8 U3927 ( .A(n2527), .B(n2232), .Z(n2257) );
  ND2SVTX4 U3928 ( .A(n1756), .B(n892), .Z(n2258) );
  ND3ASVTX8 U3929 ( .A(n2742), .B(n2260), .C(n3240), .Z(n3654) );
  IVSVTX4 U3930 ( .A(n2892), .Z(n2261) );
  ND2SVTX8 U3931 ( .A(n2741), .B(n2263), .Z(n3673) );
  ND2SVTX4 U3932 ( .A(n733), .B(n3378), .Z(n2267) );
  AO6SVTX8 U3933 ( .A(n4260), .B(n4258), .C(n2367), .Z(n4248) );
  AO7SVTX8 U3934 ( .A(n2281), .B(n2280), .C(n2546), .Z(n2282) );
  ND2SVTX6 U3935 ( .A(n2529), .B(n2531), .Z(n2280) );
  ND2SVTX6 U3936 ( .A(n3588), .B(n3589), .Z(n3593) );
  ND3SVTX4 U3937 ( .A(n575), .B(n793), .C(n4024), .Z(n4027) );
  CTIVSVTX4 U3938 ( .A(n623), .Z(n2285) );
  NR2ASVTX6 U3939 ( .A(n1112), .B(n2287), .Z(n2558) );
  ND2SVTX4 U3940 ( .A(n2305), .B(n2307), .Z(n2707) );
  ND2SVTX4 U3941 ( .A(n2290), .B(n3122), .Z(n3148) );
  NR2SVTX4 U3942 ( .A(n3970), .B(n3686), .Z(n2296) );
  ND2SVTX4 U3943 ( .A(n2295), .B(n2620), .Z(n2571) );
  IVSVTX4 U3944 ( .A(n2540), .Z(n2295) );
  IVSVTX4 U3945 ( .A(n2681), .Z(n2611) );
  ND2SVTX4 U3946 ( .A(n2583), .B(n2299), .Z(n2681) );
  NR2ASVTX6 U3947 ( .A(n640), .B(n2333), .Z(n2299) );
  AN2SVTX8 U3948 ( .A(n2782), .B(n2783), .Z(n2788) );
  F_ENSVTX2 U3949 ( .A(n3891), .B(n3890), .Z(n2315) );
  NR2SVTX4 U3950 ( .A(num_i[23]), .B(num_i[22]), .Z(n2498) );
  ND2SVTX6 U3951 ( .A(n3594), .B(n2402), .Z(n2324) );
  F_ENSVTX2 U3952 ( .A(n622), .B(n615), .Z(n2328) );
  ND2SVTX4 U3953 ( .A(n2338), .B(n2455), .Z(n3848) );
  IVSVTX4 U3954 ( .A(n2337), .Z(n2455) );
  NR2SVTX2 U3955 ( .A(n2370), .B(n1339), .Z(n2896) );
  NR2SVTX2 U3956 ( .A(n697), .B(n3536), .Z(n3537) );
  IVSVTX2 U3957 ( .A(n3214), .Z(n2345) );
  ND2SVTX4 U3958 ( .A(n4110), .B(n961), .Z(n3145) );
  IVSVTX8 U3959 ( .A(n523), .Z(n2349) );
  AO7ASVTX6 U3960 ( .A(n3768), .B(n3767), .C(n2405), .Z(n3770) );
  AO7ABSVTX8 U3961 ( .A(n2513), .B(n2126), .C(n2562), .Z(n2651) );
  ND2SVTX2 U3962 ( .A(n3565), .B(n3564), .Z(n3576) );
  ND2SVTX4 U3963 ( .A(n2373), .B(n1665), .Z(n2354) );
  ENSVTX4 U3964 ( .A(n4276), .B(n4275), .Z(rslt_o[21]) );
  IVSVTX2 U3965 ( .A(n3557), .Z(n3474) );
  NR2ASVTX2 U3966 ( .A(n3270), .B(n765), .Z(n3380) );
  NR2ASVTX2 U3967 ( .A(n3502), .B(n3501), .Z(n3507) );
  AO7NSVTX4 U3968 ( .A(n697), .B(n4020), .C(n4019), .Z(n2445) );
  ND2SVTX4 U3969 ( .A(n1688), .B(n429), .Z(n4259) );
  ND2SVTX4 U3970 ( .A(n3813), .B(n3093), .Z(n3823) );
  ND3SVTX2 U3971 ( .A(n3111), .B(n3054), .C(n3053), .Z(n3047) );
  ND4SVTX6 U3972 ( .A(n3646), .B(n3648), .C(n3649), .D(n3647), .Z(n3650) );
  AO17SVTX4 U3973 ( .A(n3633), .B(n2401), .C(n2458), .D(n3613), .Z(n3649) );
  IVSVTX2 U3974 ( .A(n3796), .Z(n2363) );
  ND2ASVTX1 U3975 ( .A(n553), .B(n2582), .Z(n2583) );
  ND3SVTX4 U3976 ( .A(n1883), .B(n3771), .C(n3986), .Z(n3776) );
  F_EOSVTX2 U3977 ( .A(n2344), .B(n606), .Z(n3035) );
  AO7ABSVTX4 U3978 ( .A(n2796), .B(n591), .C(n2417), .Z(n2797) );
  AO6SVTX2 U3979 ( .A(n4014), .B(n3939), .C(n4009), .Z(n3785) );
  NR4ABCSVTX8 U3980 ( .A(n508), .B(n545), .C(n643), .D(n2642), .Z(n2724) );
  NR3SVTX2 U3981 ( .A(n4000), .B(n4001), .C(n1697), .Z(n4002) );
  IVSVTX2 U3982 ( .A(n4290), .Z(n4191) );
  AO7SVTX2 U3983 ( .A(n3653), .B(n3655), .C(n3568), .Z(n3578) );
  AO7ASVTX2 U3984 ( .A(n2427), .B(n1690), .C(n3599), .Z(n3600) );
  NR2SVTX2 U3985 ( .A(n1791), .B(n3272), .Z(n3384) );
  IVSVTX2 U3986 ( .A(n944), .Z(n3272) );
  AO5NSVTX2 U3987 ( .A(n2784), .B(n1759), .C(n1346), .Z(n2392) );
  FAS1SVTX4 U3988 ( .A(n2348), .B(n3270), .CI(n1254), .CO(n2923), .Z(n2921) );
  IVSVTX2 U3989 ( .A(n3664), .Z(n3680) );
  IVSVTX8 U3990 ( .A(n1025), .Z(n2887) );
  AO7ABSVTX4 U3991 ( .A(n2887), .B(n2986), .C(n2985), .Z(n2987) );
  F_AN2SVTX2 U3992 ( .A(n3543), .B(n3544), .Z(n2450) );
  NR2SVTX2 U3993 ( .A(n2149), .B(n765), .Z(n3892) );
  F_ND2ASVTX2 U3994 ( .A(n3281), .B(n3642), .Z(n3643) );
  F_ENSVTX2 U3995 ( .A(n3507), .B(n3506), .Z(n3514) );
  IVSVTX2 U3996 ( .A(n4127), .Z(n4128) );
  ND2SVTX4 U3997 ( .A(n2868), .B(n2791), .Z(n2793) );
  NR2SVTX2 U3998 ( .A(n4296), .B(n1720), .Z(n4300) );
  IVSVTX4 U3999 ( .A(n799), .Z(n3509) );
  ND2SVTX4 U4000 ( .A(n1596), .B(n3799), .Z(n3800) );
  NR2SVTX2 U4001 ( .A(n1347), .B(n942), .Z(n4005) );
  AO6CSVTX6 U4002 ( .A(n1744), .B(n2524), .C(n2523), .Z(n2546) );
  IVSVTX2 U4003 ( .A(n3401), .Z(n3404) );
  ND2ASVTX8 U4004 ( .A(n2589), .B(n2552), .Z(n2539) );
  BFSVTX4 U4005 ( .A(num_i[29]), .Z(n2695) );
  AO7SVTX2 U4006 ( .A(n652), .B(n3122), .C(n1741), .Z(n2870) );
  NR2ASVTX2 U4007 ( .A(n4171), .B(n4021), .Z(n4028) );
  AN2SVTX4 U4008 ( .A(n445), .B(n2009), .Z(n2425) );
  IVSVTX2 U4009 ( .A(n3138), .Z(n2869) );
  F_ND2ASVTX2 U4010 ( .A(n2760), .B(n3078), .Z(n2761) );
  IVSVTX2 U4011 ( .A(n3594), .Z(n3541) );
  ND3ASVTX2 U4012 ( .A(n3543), .B(n3594), .C(n3540), .Z(n3549) );
  AO7ABSVTX2 U4013 ( .A(n741), .B(n3341), .C(n3387), .Z(n3293) );
  AO7SVTX4 U4014 ( .A(n4036), .B(n4034), .C(n4035), .Z(n4040) );
  IVSVTX2 U4015 ( .A(n3006), .Z(n2966) );
  F_AN2SVTX2 U4016 ( .A(n3166), .B(n3165), .Z(n3188) );
  IVSVTX2 U4017 ( .A(n3573), .Z(n3437) );
  AO1ASVTX4 U4018 ( .A(n3111), .B(n775), .C(n573), .D(n4132), .Z(n4134) );
  IVSVTX2 U4019 ( .A(n3450), .Z(n2745) );
  IVSVTX2 U4020 ( .A(n2762), .Z(n2764) );
  F_ENSVTX2 U4021 ( .A(n3553), .B(n3512), .Z(n3513) );
  AO7SVTX4 U4022 ( .A(n3554), .B(n3553), .C(n799), .Z(n3555) );
  ND3SVTX4 U4023 ( .A(n3822), .B(n3823), .C(n3821), .Z(n3826) );
  CTIVSVTX2 U4024 ( .A(n3774), .Z(n3769) );
  IVSVTX4 U4025 ( .A(n3798), .Z(n3801) );
  NR2SVTX2 U4026 ( .A(n3191), .B(n3168), .Z(n3169) );
  ND2SVTX4 U4027 ( .A(n3635), .B(n2401), .Z(n3647) );
  IVSVTX2 U4028 ( .A(n2354), .Z(n3627) );
  NR2SVTX2 U4029 ( .A(n3576), .B(n3574), .Z(n3575) );
  AO7SVTX2 U4030 ( .A(n3576), .B(n3569), .C(n2424), .Z(n3581) );
  IVSVTX2 U4031 ( .A(n3578), .Z(n3569) );
  ND2SVTX2 U4032 ( .A(n3260), .B(n523), .Z(n3269) );
  AO7CSVTX4 U4033 ( .A(n4082), .B(n4081), .C(n4080), .Z(n4083) );
  AO7SVTX2 U4034 ( .A(n4079), .B(n571), .C(n1596), .Z(n4080) );
  IVSVTX2 U4035 ( .A(n2685), .Z(n2691) );
  IVSVTX2 U4036 ( .A(n3834), .Z(n3832) );
  NR2SVTX2 U4037 ( .A(n3897), .B(n3895), .Z(n3894) );
  IVSVTX2 U4038 ( .A(n3852), .Z(n3766) );
  AO7SVTX2 U4039 ( .A(n3533), .B(n3534), .C(n3532), .Z(n3479) );
  IVSVTX2 U4040 ( .A(n3952), .Z(n3953) );
  IVSVTX2 U4041 ( .A(n3244), .Z(n3173) );
  AO2ABSVTX4 U4042 ( .C(n3192), .D(n3168), .A(n3191), .B(n1270), .Z(n3193) );
  IVSVTX2 U4043 ( .A(n3028), .Z(n3124) );
  IVSVTX2 U4044 ( .A(n3658), .Z(n3657) );
  IVSVTX2 U4045 ( .A(n3712), .Z(n3705) );
  F_ND2ASVTX2 U4046 ( .A(n3949), .B(n1422), .Z(n3934) );
  IVSVTX2 U4047 ( .A(n3409), .Z(n3410) );
  F_MUX21NSVTX1 U4048 ( .A(n3359), .B(n3384), .S(n3362), .Z(n3360) );
  B_ND2SVTX2 U4049 ( .A(n2465), .B(n3363), .Z(n3364) );
  AO3SVTX2 U4050 ( .A(n3307), .B(n3366), .C(n3306), .D(n4066), .Z(n3308) );
  NR2SVTX2 U4051 ( .A(n2248), .B(n4043), .Z(n4044) );
  F_ND2ASVTX2 U4052 ( .A(n4033), .B(n4032), .Z(n4046) );
  NR2SVTX2 U4053 ( .A(n4041), .B(n4039), .Z(n4033) );
  F_ND3SVTX2 U4054 ( .A(n4174), .B(n367), .C(n4173), .Z(n4182) );
  AO7SVTX2 U4055 ( .A(n4197), .B(n1678), .C(n4148), .Z(n4087) );
  AO7ABSVTX4 U4056 ( .A(n592), .B(n3857), .C(n3854), .Z(n3864) );
  ND3SVTX4 U4057 ( .A(n3576), .B(n3568), .C(n3574), .Z(n3567) );
  ND3SVTX4 U4058 ( .A(n2644), .B(n1805), .C(n2126), .Z(n2645) );
  IVSVTX4 U4059 ( .A(n3101), .Z(n3104) );
  IVSVTX2 U4060 ( .A(n3787), .Z(n3743) );
  NR2ASVTX2 U4061 ( .A(n4160), .B(n560), .Z(n4155) );
  NR2ASVTX2 U4062 ( .A(n2698), .B(n1544), .Z(n2630) );
  NR2ASVTX2 U4063 ( .A(n2369), .B(n2561), .Z(n2553) );
  F_ND2SVTX0H U4064 ( .A(n4190), .B(n4189), .Z(n4193) );
  ND2SVTX2 U4065 ( .A(n1789), .B(n3272), .Z(n3386) );
  FAS1SVTX4 U4066 ( .A(n1419), .B(n2812), .CI(n944), .CO(n2818), .Z(n2816) );
  AO5ASVTX6 U4067 ( .B(n508), .A(n2888), .C(n2887), .Z(n2889) );
  IVSVTX0H U4068 ( .A(n4248), .Z(n4256) );
  IVSVTX2 U4069 ( .A(n3382), .Z(n3353) );
  ND2SVTX2 U4070 ( .A(n570), .B(n3382), .Z(n3409) );
  ND2ASVTX8 U4071 ( .A(n3456), .B(n3455), .Z(n3473) );
  ND2SVTX4 U4072 ( .A(n3074), .B(n3073), .Z(n3453) );
  F_ND2ASVTX2 U4073 ( .A(n540), .B(n3126), .Z(n2956) );
  F_EOSVTX2 U4074 ( .A(n2344), .B(n622), .Z(n2941) );
  NR2ASVTX1 U4075 ( .A(n4176), .B(n4175), .Z(n4177) );
  ND3ABSVTX4 U4076 ( .A(n3206), .B(n1635), .C(n2139), .Z(n3209) );
  IVSVTX2 U4077 ( .A(n2854), .Z(n2855) );
  NR2SVTX4 U4078 ( .A(n3632), .B(n3631), .Z(n2401) );
  AO2SVTX4 U4079 ( .A(n3752), .B(n3753), .C(n3751), .D(n2397), .Z(n3756) );
  ND3ABSVTX4 U4080 ( .A(n2397), .B(n3749), .C(n2463), .Z(n3750) );
  F_AN2SVTX2 U4081 ( .A(n3748), .B(n3747), .Z(n2397) );
  F_EOSVTX2 U4082 ( .A(n3126), .B(n3014), .Z(n2927) );
  ND2SVTX4 U4083 ( .A(n2167), .B(n4124), .Z(n4125) );
  AO5SVTX2 U4084 ( .A(n3014), .B(n2720), .C(n2392), .Z(n3025) );
  IVSVTX2 U4085 ( .A(n3701), .Z(n3716) );
  IVSVTX6 U4086 ( .A(n878), .Z(n3613) );
  F_EOSVTX2 U4087 ( .A(n1642), .B(n2776), .Z(n2794) );
  AO7SVTX6 U4088 ( .A(n1932), .B(n3051), .C(n459), .Z(n3097) );
  ND2SVTX4 U4089 ( .A(n3737), .B(n3738), .Z(n3740) );
  NR2ASVTX2 U4090 ( .A(n2940), .B(n3342), .Z(n3345) );
  IVSVTX2 U4091 ( .A(n413), .Z(n4289) );
  NR2SVTX2 U4092 ( .A(n2344), .B(n2743), .Z(n2388) );
  ND2SVTX4 U4093 ( .A(n3332), .B(n3170), .Z(n3336) );
  AO7SVTX4 U4094 ( .A(n775), .B(n3126), .C(n1494), .Z(n4074) );
  AO3SVTX4 U4095 ( .A(n3068), .B(n1089), .C(n1397), .D(n814), .Z(n2734) );
  NR2SVTX2 U4096 ( .A(n2611), .B(n2898), .Z(n2694) );
  AN2SVTX4 U4097 ( .A(n891), .B(n513), .Z(n2409) );
  AO7SVTX4 U4098 ( .A(n3100), .B(n2971), .C(n3099), .Z(n3101) );
  AO7SVTX4 U4099 ( .A(n895), .B(n2578), .C(n1629), .Z(n2581) );
  EOSVTX4 U4100 ( .A(n4253), .B(n4252), .Z(rslt_o[5]) );
  AO6SVTX2 U4101 ( .A(n4256), .B(n4249), .C(n4251), .Z(n4252) );
  ND2SVTX4 U4102 ( .A(n514), .B(n3259), .Z(n3261) );
  NR2ASVTX2 U4103 ( .A(n3920), .B(n3914), .Z(n3915) );
  IVSVTX4 U4104 ( .A(n3918), .Z(n3914) );
  ND2SVTX4 U4105 ( .A(n3911), .B(n2457), .Z(n3918) );
  IVSVTX2 U4106 ( .A(n2389), .Z(n2488) );
  ND2SVTX4 U4107 ( .A(n3460), .B(n3459), .Z(n3557) );
  ND2SVTX4 U4108 ( .A(n2385), .B(n2964), .Z(n3322) );
  FAS1SVTX4 U4109 ( .A(n3032), .B(n2789), .CI(n1642), .CO(n2787), .Z(n2799) );
  IVSVTX2 U4110 ( .A(n4221), .Z(n4279) );
  AO7ABSVTX2 U4111 ( .A(n2887), .B(n2764), .C(n2763), .Z(n2765) );
  BFSVTX12 U4112 ( .A(n4138), .Z(n4066) );
  ND2SVTX4 U4113 ( .A(n865), .B(n4086), .Z(n4148) );
  AN2SVTX4 U4114 ( .A(n3748), .B(n3784), .Z(n2416) );
  NR2ASVTX6 U4115 ( .A(n3111), .B(n3037), .Z(n3247) );
  F_IVSVTX0H U4116 ( .A(num_i[6]), .Z(n2631) );
  F_IVSVTX0H U4117 ( .A(n3808), .Z(n3610) );
  ENSVTX0H U4118 ( .A(n3286), .B(n2747), .Z(n2454) );
  NR3SVTX2 U4119 ( .A(num_i[16]), .B(n2584), .C(n2573), .Z(n2490) );
  F_AN2SVTX2 U4120 ( .A(n3222), .B(n4055), .Z(n2461) );
  AN2SVTX0H U4121 ( .A(n3362), .B(n3386), .Z(n2465) );
  IVSVTX4 U4122 ( .A(n1591), .Z(n4069) );
  IVSVTX4 U4123 ( .A(n545), .Z(n3078) );
  NR2SVTX4 U4124 ( .A(num_i[5]), .B(num_i[4]), .Z(n2469) );
  AO7SVTX4 U4125 ( .A(num_i[2]), .B(num_i[3]), .C(n2469), .Z(n2471) );
  ND2SVTX4 U4126 ( .A(n2471), .B(n2470), .Z(n2477) );
  NR2SVTX8 U4127 ( .A(num_i[20]), .B(num_i[21]), .Z(n2497) );
  IVSVTX4 U4128 ( .A(num_i[23]), .Z(n2478) );
  IVSVTX4 U4129 ( .A(num_i[22]), .Z(n2518) );
  BFSVTX12 U4130 ( .A(num_i[18]), .Z(n2584) );
  NR2SVTX4 U4131 ( .A(num_i[17]), .B(num_i[24]), .Z(n2492) );
  NR2SVTX6 U4132 ( .A(num_i[31]), .B(num_i[17]), .Z(n2500) );
  IVSVTX4 U4133 ( .A(num_i[5]), .Z(n2646) );
  NR2SVTX2 U4134 ( .A(num_i[6]), .B(n2646), .Z(n2510) );
  NR2ASVTX6 U4135 ( .A(n2577), .B(n2522), .Z(n2524) );
  IVSVTX4 U4136 ( .A(num_i[30]), .Z(n2682) );
  AO6SVTX2 U4137 ( .A(n2682), .B(num_i[29]), .C(num_i[31]), .Z(n2523) );
  NR2SVTX8 U4138 ( .A(n2533), .B(n2532), .Z(n2657) );
  CTBUFSVTX2 U4139 ( .A(num_i[12]), .Z(n2579) );
  ND2SVTX4 U4140 ( .A(n2539), .B(n2538), .Z(n2623) );
  IVSVTX0H U4141 ( .A(n2573), .Z(n2574) );
  ND2SVTX6 U4142 ( .A(n2595), .B(n2594), .Z(n2609) );
  ND2SVTX8 U4143 ( .A(n2604), .B(n2603), .Z(n2947) );
  AO7SVTX2 U4144 ( .A(n2518), .B(n895), .C(n2682), .Z(n2690) );
  IVSVTX2 U4145 ( .A(n2690), .Z(n2684) );
  AN2SVTX8 U4146 ( .A(n2701), .B(n2702), .Z(n2720) );
  ND3SVTX4 U4147 ( .A(n1686), .B(n546), .C(n2734), .Z(n2739) );
  IVSVTX4 U4148 ( .A(n2882), .Z(n3452) );
  ND2SVTX4 U4149 ( .A(n428), .B(n2883), .Z(n3450) );
  IVSVTX2 U4150 ( .A(n3440), .Z(n2754) );
  ND2SVTX2 U4151 ( .A(n3079), .B(n2758), .Z(n3073) );
  NR2ASVTX6 U4152 ( .A(n2769), .B(n2768), .Z(rslt_o[0]) );
  AO5SVTX4 U4153 ( .A(n444), .B(n2788), .C(n621), .Z(n2798) );
  NR2ASVTX8 U4154 ( .A(n2804), .B(n2803), .Z(n3211) );
  ND3SVTX8 U4155 ( .A(n2837), .B(n2836), .C(n3668), .Z(n2843) );
  ND3SVTX8 U4156 ( .A(n3620), .B(n3619), .C(n3618), .Z(n2860) );
  IVSVTX2 U4157 ( .A(n2846), .Z(n2847) );
  NR2SVTX4 U4158 ( .A(n2412), .B(n2928), .Z(n3138) );
  IVSVTX2 U4159 ( .A(n2922), .Z(n2872) );
  FAS1SVTX4 U4160 ( .A(n709), .B(n1025), .CI(n2905), .CO(n2878), .Z(n2881) );
  NR2SVTX4 U4161 ( .A(n517), .B(n2316), .Z(n2886) );
  NR2SVTX8 U4162 ( .A(n2889), .B(n2890), .Z(n3554) );
  FAS1SVTX4 U4163 ( .A(n1361), .B(n1881), .CI(n2993), .CO(n2916), .Z(n2914) );
  AO7SVTX2 U4164 ( .A(n3166), .B(n3138), .C(n3137), .Z(n4101) );
  IVSVTX2 U4165 ( .A(n3035), .Z(n3034) );
  NR2ASVTX2 U4166 ( .A(n2931), .B(n3034), .Z(n4145) );
  ND2SVTX4 U4167 ( .A(n2953), .B(n2952), .Z(n3201) );
  ND2SVTX4 U4168 ( .A(n2956), .B(n1789), .Z(n2957) );
  ND2SVTX4 U4169 ( .A(n2966), .B(n2965), .Z(n3956) );
  FAS1SVTX4 U4170 ( .A(n1295), .B(n2971), .CI(n1743), .CO(n3006), .Z(n3723) );
  ND2SVTX8 U4171 ( .A(n600), .B(n3004), .Z(n3722) );
  ND2SVTX4 U4172 ( .A(n605), .B(n2999), .Z(n3591) );
  IVSVTX0H U4173 ( .A(n4147), .Z(n3110) );
  FAS1SVTX4 U4174 ( .A(n3311), .B(n2344), .CI(n3022), .CO(n3027), .Z(n3037) );
  CTIVSVTX4 U4175 ( .A(n3027), .Z(n3023) );
  ND2SVTX8 U4176 ( .A(n1923), .B(n3023), .Z(n3244) );
  NR3ABSVTX8 U4177 ( .A(n3244), .B(n3028), .C(n3026), .Z(n4151) );
  ND2SVTX2 U4178 ( .A(n3039), .B(n3040), .Z(n3312) );
  ND2ASVTX8 U4179 ( .A(n3060), .B(n3089), .Z(n3818) );
  NR2SVTX8 U4180 ( .A(n3082), .B(n3081), .Z(n3501) );
  ND2SVTX4 U4181 ( .A(n3082), .B(n3081), .Z(n3502) );
  ND2SVTX4 U4182 ( .A(n3094), .B(n3095), .Z(n3871) );
  IVSVTX4 U4183 ( .A(n3098), .Z(n3100) );
  ND2SVTX6 U4184 ( .A(n3104), .B(n3103), .Z(n3787) );
  ND2SVTX4 U4185 ( .A(n3175), .B(n3244), .Z(n3129) );
  AO7SVTX4 U4186 ( .A(n3127), .B(n3245), .C(n3174), .Z(n3128) );
  ND2SVTX4 U4187 ( .A(n3136), .B(n3134), .Z(n3130) );
  ND2SVTX4 U4188 ( .A(n3131), .B(n3130), .Z(n3133) );
  IVSVTX4 U4189 ( .A(n3142), .Z(n3168) );
  IVSVTX0H U4190 ( .A(n3166), .Z(n3140) );
  IVSVTX2 U4191 ( .A(n3151), .Z(n3202) );
  ND2SVTX4 U4192 ( .A(n2393), .B(n2009), .Z(n4132) );
  IVSVTX4 U4193 ( .A(n4132), .Z(n3160) );
  ND2ASVTX8 U4194 ( .A(n3161), .B(n3160), .Z(n4075) );
  ND2SVTX2 U4195 ( .A(n4138), .B(n3167), .Z(n3191) );
  IVSVTX4 U4196 ( .A(n4032), .Z(n4037) );
  ND2SVTX4 U4197 ( .A(n3175), .B(n3174), .Z(n3180) );
  AO6SVTX4 U4198 ( .A(n3179), .B(n3178), .C(n3177), .Z(n3182) );
  ND2SVTX2 U4199 ( .A(n3217), .B(n3216), .Z(n3218) );
  NR3ABSVTX4 U4200 ( .A(n3351), .B(n3220), .C(n573), .Z(n3257) );
  ND3SVTX2 U4201 ( .A(n3235), .B(n3236), .C(n3237), .Z(n3238) );
  ND3SVTX2 U4202 ( .A(n2461), .B(n3239), .C(n3238), .Z(n3243) );
  ND2SVTX2 U4203 ( .A(n3245), .B(n3244), .Z(n3254) );
  AO7SVTX4 U4204 ( .A(n3248), .B(n3333), .C(n3170), .Z(n3253) );
  NR2SVTX4 U4205 ( .A(n3254), .B(n3253), .Z(n3250) );
  AO7SVTX2 U4206 ( .A(n3254), .B(n3332), .C(n1422), .Z(n3249) );
  NR2SVTX4 U4207 ( .A(n3261), .B(n2361), .Z(n3263) );
  F_AN2SVTX2 U4208 ( .A(n3267), .B(n3323), .Z(n3268) );
  NR2SVTX2 U4209 ( .A(n1743), .B(n3270), .Z(n3356) );
  NR2SVTX2 U4210 ( .A(n3384), .B(n3356), .Z(n3341) );
  AO7SVTX4 U4211 ( .A(n3356), .B(n3386), .C(n3358), .Z(n3342) );
  AO7SVTX6 U4212 ( .A(n3532), .B(n614), .C(n3478), .Z(n3675) );
  ND2SVTX4 U4213 ( .A(n964), .B(n1033), .Z(n3495) );
  AO6SVTX4 U4214 ( .A(n3749), .B(n3748), .C(n3746), .Z(n4006) );
  IVSVTX0H U4215 ( .A(n3366), .Z(n3302) );
  ND3SVTX8 U4216 ( .A(n533), .B(n482), .C(n1321), .Z(n3369) );
  F_ND2ASVTX2 U4217 ( .A(n3311), .B(n3310), .Z(n3365) );
  NR2SVTX4 U4218 ( .A(n3315), .B(n3313), .Z(n3314) );
  AO17SVTX2 U4219 ( .A(n3341), .B(n741), .C(n2385), .D(n1609), .Z(n3346) );
  ND2SVTX4 U4220 ( .A(n3352), .B(n3351), .Z(n3355) );
  IVSVTX2 U4221 ( .A(n3356), .Z(n3357) );
  ND2SVTX2 U4222 ( .A(n3358), .B(n3357), .Z(n3362) );
  ND2SVTX4 U4223 ( .A(n3370), .B(n3371), .Z(n3379) );
  IVSVTX0H U4224 ( .A(n3384), .Z(n3385) );
  ND2SVTX4 U4225 ( .A(n1321), .B(n3390), .Z(n3401) );
  IVSVTX4 U4226 ( .A(n3392), .Z(n4036) );
  AO7SVTX4 U4227 ( .A(n4036), .B(n3398), .C(n3395), .Z(n3407) );
  IVSVTX4 U4228 ( .A(n3420), .Z(n3421) );
  NR2SVTX6 U4229 ( .A(n4281), .B(n4284), .Z(n4290) );
  ND2ASVTX8 U4230 ( .A(n4171), .B(n3972), .Z(n3905) );
  ND2SVTX4 U4231 ( .A(n3428), .B(n3591), .Z(n3429) );
  ND2SVTX4 U4232 ( .A(n3437), .B(n3438), .Z(n3448) );
  IVSVTX2 U4233 ( .A(n3463), .Z(n3464) );
  F_ENSVTX2 U4234 ( .A(n3480), .B(n3479), .Z(n3481) );
  ND2SVTX4 U4235 ( .A(n3485), .B(n574), .Z(n3486) );
  NR2SVTX2 U4236 ( .A(n505), .B(n3487), .Z(n3488) );
  IVSVTX4 U4237 ( .A(n3561), .Z(n3492) );
  AO6SVTX2 U4238 ( .A(n3516), .B(n3518), .C(n3515), .Z(n3496) );
  AO6CSVTX8 U4239 ( .A(n3519), .B(n3521), .C(n3508), .Z(n3553) );
  AO7SVTX8 U4240 ( .A(n3563), .B(n4248), .C(n3562), .Z(n4231) );
  ND2SVTX4 U4241 ( .A(n3656), .B(n1474), .Z(n3574) );
  NR2SVTX8 U4242 ( .A(n3593), .B(n3592), .Z(n3595) );
  ND2SVTX6 U4243 ( .A(n3594), .B(n3595), .Z(n3628) );
  ND2SVTX4 U4244 ( .A(n3809), .B(n3817), .Z(n3612) );
  NR2SVTX2 U4245 ( .A(n3624), .B(n2997), .Z(n3693) );
  ND2SVTX4 U4246 ( .A(n2373), .B(n1665), .Z(n3694) );
  ND2SVTX4 U4247 ( .A(n3808), .B(n3809), .Z(n3873) );
  IVSVTX0H U4248 ( .A(n3636), .Z(n3637) );
  NR2ASVTX1 U4249 ( .A(n3638), .B(n3637), .Z(n3644) );
  F_ENSVTX2 U4250 ( .A(n3644), .B(n3643), .Z(n3645) );
  ND2SVTX4 U4251 ( .A(n530), .B(n3645), .Z(n3646) );
  IVSVTX0H U4252 ( .A(n3675), .Z(n3670) );
  AO1SVTX4 U4253 ( .A(n3679), .B(n3675), .C(n3674), .D(n697), .Z(n3676) );
  NR2SVTX4 U4254 ( .A(n4234), .B(n3687), .Z(n3718) );
  AO7SVTX4 U4255 ( .A(n3684), .B(n2997), .C(n3691), .Z(n3695) );
  AO6SVTX8 U4256 ( .A(n4231), .B(n3718), .C(n3717), .Z(n4214) );
  ND2ASVTX8 U4257 ( .A(n1697), .B(n3928), .Z(n3727) );
  IVSVTX4 U4258 ( .A(n3924), .Z(n3720) );
  NR2SVTX8 U4259 ( .A(n4000), .B(n3720), .Z(n3726) );
  F_AN2SVTX2 U4260 ( .A(n3724), .B(n3723), .Z(n3970) );
  IVSVTX2 U4261 ( .A(n3970), .Z(n3725) );
  ND3ABSVTX8 U4262 ( .A(n3743), .B(n3740), .C(n3742), .Z(n3744) );
  NR2ASVTX2 U4263 ( .A(n3852), .B(n3856), .Z(n3774) );
  IVSVTX0H U4264 ( .A(n3893), .Z(n3768) );
  F_ND2SVTX0H U4265 ( .A(n3784), .B(n3783), .Z(n3786) );
  ND2SVTX4 U4266 ( .A(n3802), .B(n3928), .Z(n3799) );
  ND2SVTX6 U4267 ( .A(n3805), .B(n3804), .Z(n3806) );
  IVSVTX4 U4268 ( .A(n3814), .Z(n3932) );
  CTIVSVTX4 U4269 ( .A(n3932), .Z(n3820) );
  NR2ASVTX6 U4270 ( .A(n3818), .B(n2452), .Z(n3879) );
  AO7ABSVTX6 U4271 ( .A(n3820), .B(n3930), .C(n3819), .Z(n3821) );
  NR2SVTX8 U4272 ( .A(n3828), .B(n602), .Z(n3835) );
  NR2ASVTX6 U4273 ( .A(n3886), .B(n3835), .Z(n3834) );
  ND2SVTX2 U4274 ( .A(n3834), .B(n926), .Z(n3837) );
  ND3SVTX2 U4275 ( .A(n3887), .B(n3835), .C(n3889), .Z(n3836) );
  NR2ASVTX2 U4276 ( .A(n3858), .B(n3857), .Z(n3860) );
  ND2SVTX4 U4277 ( .A(n3860), .B(n3859), .Z(n3861) );
  ND2SVTX4 U4278 ( .A(n3896), .B(n3986), .Z(n3901) );
  NR2SVTX2 U4279 ( .A(n569), .B(n587), .Z(n3913) );
  IVSVTX4 U4280 ( .A(n2200), .Z(n3925) );
  F_AN2SVTX2 U4281 ( .A(n4035), .B(n415), .Z(n3949) );
  NR3SVTX2 U4282 ( .A(n3939), .B(n3938), .C(n3937), .Z(n3943) );
  NR3SVTX2 U4283 ( .A(n4011), .B(n3945), .C(n3941), .Z(n3942) );
  IVSVTX2 U4284 ( .A(n3974), .Z(n3976) );
  IVSVTX2 U4285 ( .A(n1409), .Z(n3997) );
  AO6SVTX2 U4286 ( .A(n4009), .B(n4010), .C(n4008), .Z(n4015) );
  NR2SVTX4 U4287 ( .A(n4012), .B(n4011), .Z(n4013) );
  F_ENSVTX2 U4288 ( .A(n4017), .B(n4016), .Z(n4020) );
  MUX21NSVTX2 U4289 ( .A(n4042), .B(n4041), .S(n4040), .Z(n4043) );
  ND2SVTX6 U4290 ( .A(n4220), .B(n4052), .Z(n4053) );
  NR3SVTX4 U4291 ( .A(n4063), .B(n4062), .C(n4061), .Z(n4064) );
  AO7SVTX2 U4292 ( .A(n2385), .B(n4069), .C(n4068), .Z(n4072) );
  AO6ABSVTX4 U4293 ( .A(n2940), .B(n1591), .C(n4070), .Z(n4071) );
  EOSVTX8 U4294 ( .A(n4090), .B(n4089), .Z(rslt_o[22]) );
  NR2SVTX2 U4295 ( .A(n4145), .B(n1983), .Z(n4102) );
  IVSVTX4 U4296 ( .A(n4122), .Z(n4178) );
  IVSVTX2 U4297 ( .A(n4123), .Z(n4124) );
  F_AN2SVTX2 U4298 ( .A(n4163), .B(n3854), .Z(n4142) );
  AO20SVTX2 U4299 ( .A(n4158), .B(n4157), .C(n4163), .D(n2248), .Z(n4161) );
  AO2SVTX2 U4300 ( .A(n4167), .B(n4168), .C(n2349), .D(n367), .Z(n4170) );
  AO20SVTX2 U4301 ( .A(n2167), .B(n4178), .C(n4177), .D(n2776), .Z(n4181) );
  AO7ABSVTX4 U4302 ( .A(n2440), .B(n4185), .C(n4184), .Z(n4203) );
  ND2SVTX4 U4303 ( .A(n4206), .B(n4203), .Z(n4188) );
  NR2SVTX2 U4304 ( .A(n4191), .B(n413), .Z(n4192) );
  ND2SVTX2 U4305 ( .A(n4204), .B(n1659), .Z(n4195) );
  EOSVTX8 U4306 ( .A(n4195), .B(n4187), .Z(rslt_o[23]) );
  ND2SVTX2 U4307 ( .A(n556), .B(n4197), .Z(n4199) );
  EOSVTX8 U4308 ( .A(n4199), .B(n4198), .Z(rslt_o[20]) );
  EOSVTX8 U4309 ( .A(n4212), .B(n4211), .Z(rslt_o[25]) );
  IVSVTX2 U4310 ( .A(n4214), .Z(n4301) );
  IVSVTX0H U4311 ( .A(n4215), .Z(n4242) );
  BFSVTX1 U4312 ( .A(n4216), .Z(n4241) );
  IVSVTX2 U4313 ( .A(n4231), .Z(n4245) );
  ND2SVTX2 U4314 ( .A(n4244), .B(n4229), .Z(n4238) );
  ND2SVTX2 U4315 ( .A(n4242), .B(n4241), .Z(n4243) );
  BFSVTX1 U4316 ( .A(n4250), .Z(n4254) );
  BFSVTX1 U4317 ( .A(n4261), .Z(n4265) );
  IVSVTX2 U4318 ( .A(n1678), .Z(n4269) );
  IVSVTX0H U4319 ( .A(n4281), .Z(n4282) );
  ND2SVTX2 U4320 ( .A(n4282), .B(n4283), .Z(n4287) );
  AO6SVTX4 U4321 ( .A(n4306), .B(n4304), .C(n4285), .Z(n4286) );
  EOSVTX4 U4322 ( .A(n4287), .B(n4286), .Z(rslt_o[16]) );
  IVSVTX0H U4323 ( .A(n4295), .Z(n4296) );
  AO6SVTX2 U4324 ( .A(n4301), .B(n4300), .C(n4299), .Z(n4302) );
  EOSVTX4 U4325 ( .A(n4303), .B(n4302), .Z(rslt_o[12]) );
endmodule

