
module remap ( m1, m2 );
  input [27:0] m1;
  output [26:0] m2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664;

  F_ENSVTX2 U3 ( .A(n1384), .B(n1383), .Z(m2[16]) );
  ENSVTX6 U4 ( .A(n1345), .B(n1344), .Z(m2[21]) );
  NR2ASVTX1 U5 ( .A(n1160), .B(n985), .Z(n1165) );
  AO1SVTX1 U6 ( .A(n1296), .B(n1628), .C(n1627), .D(n1626), .Z(n1629) );
  IVSVTX0H U7 ( .A(n1317), .Z(n1307) );
  AO7SVTX1 U8 ( .A(n1238), .B(n1598), .C(n1597), .Z(n1599) );
  NR3SVTX6 U9 ( .A(n1042), .B(n990), .C(n993), .Z(n991) );
  NR4ABSVTX6 U10 ( .A(n1299), .B(n1247), .C(n1246), .D(n1245), .Z(n1259) );
  ENSVTX0H U11 ( .A(n1175), .B(n1174), .Z(n1206) );
  EOSVTX0H U12 ( .A(n1350), .B(n1349), .Z(n1380) );
  ENSVTX0H U13 ( .A(n1262), .B(n1261), .Z(n1298) );
  NR2ASVTX1 U14 ( .A(n1352), .B(n1353), .Z(n1262) );
  NR2ASVTX1 U15 ( .A(n1633), .B(n1635), .Z(n1175) );
  IVSVTX2 U16 ( .A(n1152), .Z(n1155) );
  IVSVTX0H U17 ( .A(n1300), .Z(n1301) );
  CTIVSVTX2 U18 ( .A(n1335), .Z(n1336) );
  AO7SVTX1 U19 ( .A(n1501), .B(n1503), .C(n1502), .Z(n1422) );
  AO7SVTX1 U20 ( .A(n1260), .B(n1606), .C(n441), .Z(n1261) );
  AO6NSVTX1 U21 ( .A(n1310), .B(n1309), .C(n1308), .Z(n1330) );
  NR2ASVTX1 U22 ( .A(n1589), .B(n1591), .Z(n1552) );
  IVSVTX0H U23 ( .A(n1602), .Z(n1604) );
  IVSVTX0H U24 ( .A(n1323), .Z(n1326) );
  BFSVTX4 U25 ( .A(n1163), .Z(n1335) );
  AO6SVTX1 U26 ( .A(n1644), .B(n120), .C(n119), .Z(n1349) );
  IVSVTX0H U27 ( .A(n385), .Z(n101) );
  NR2ASVTX4 U28 ( .A(n1253), .B(n1041), .Z(n989) );
  OR2SVTX2 U29 ( .A(n1242), .B(n1241), .Z(n1258) );
  BFSVTX2 U30 ( .A(n1650), .Z(n45) );
  IVSVTX0H U31 ( .A(n1460), .Z(n1497) );
  NR2ASVTX1 U32 ( .A(n1647), .B(n1646), .Z(n1656) );
  IVSVTX0H U33 ( .A(n1458), .Z(n1471) );
  IVSVTX0H U34 ( .A(n1314), .Z(n1316) );
  AO7SVTX1 U35 ( .A(n39), .B(n1239), .C(n1238), .Z(n1242) );
  IVSVTX0H U36 ( .A(n996), .Z(n1388) );
  IVSVTX0H U37 ( .A(n1260), .Z(n1356) );
  NR2ASVTX4 U38 ( .A(n1327), .B(n1163), .Z(n1244) );
  IVSVTX0H U39 ( .A(n391), .Z(n120) );
  IVSVTX0H U40 ( .A(n1421), .Z(n1501) );
  BFSVTX4 U41 ( .A(n779), .Z(n39) );
  IVSVTX0H U42 ( .A(n1177), .Z(n1395) );
  IVSVTX0H U43 ( .A(n1452), .Z(n1484) );
  AN2BSVTX2 U44 ( .A(n156), .B(n426), .Z(n1503) );
  IVSVTX0H U45 ( .A(n1648), .Z(n1271) );
  IVSVTX0H U46 ( .A(n714), .Z(n183) );
  IVSVTX0H U47 ( .A(n1550), .Z(n1585) );
  NR2SVTX2 U48 ( .A(n1133), .B(n1132), .Z(n1147) );
  IVSVTX0H U49 ( .A(n1143), .Z(n1124) );
  AO6SVTX1 U50 ( .A(n50), .B(n1403), .C(n226), .Z(n1655) );
  IVSVTX6 U51 ( .A(n988), .Z(n1042) );
  IVSVTX0H U52 ( .A(n1002), .Z(n1498) );
  B_ND2SVTX2 U53 ( .A(n59), .B(n73), .Z(n1102) );
  AO2SVTX2 U54 ( .A(n1083), .B(n1296), .C(n1082), .D(n4), .Z(n1101) );
  IVSVTX0H U55 ( .A(n1478), .Z(n1023) );
  AO4ABSVTX4 U56 ( .C(n1123), .D(n384), .A(n1122), .B(n60), .Z(n1132) );
  AN4SVTX1 U57 ( .A(n1121), .B(n1120), .C(n26), .D(n1118), .Z(n60) );
  IVSVTX0H U58 ( .A(n1569), .Z(n150) );
  CTIVSVTX2 U59 ( .A(n941), .Z(n665) );
  IVSVTX0H U60 ( .A(n330), .Z(n50) );
  IVSVTX0H U61 ( .A(n428), .Z(n151) );
  IVSVTX0H U62 ( .A(n1025), .Z(n1027) );
  ENSVTX1 U63 ( .A(m1[24]), .B(n1074), .Z(n1083) );
  ND3ASVTX6 U64 ( .A(n806), .B(n805), .C(n804), .Z(n807) );
  AO21SVTX1 U65 ( .A(n1128), .B(n1127), .C(n1126), .D(n1061), .Z(n1129) );
  AO7SVTX2 U66 ( .A(n1057), .B(n1056), .C(n1138), .Z(n1058) );
  CTIVSVTX2 U67 ( .A(n1077), .Z(n1096) );
  ND3SVTX2 U68 ( .A(n1650), .B(n662), .C(n61), .Z(n1045) );
  IVSVTX0H U69 ( .A(n1057), .Z(n1054) );
  IVSVTX0H U70 ( .A(n1120), .Z(n1086) );
  IVSVTX0H U71 ( .A(n1012), .Z(n1013) );
  ND3ABSVTX2 U72 ( .A(n65), .B(n818), .C(n817), .Z(n1323) );
  NR2SVTX2 U73 ( .A(n778), .B(n777), .Z(n709) );
  IVSVTX0H U74 ( .A(n1121), .Z(n1091) );
  B_ND2SVTX2 U75 ( .A(n873), .B(n916), .Z(n1310) );
  ND3SVTX2 U76 ( .A(n1491), .B(n863), .C(n862), .Z(n875) );
  NR4ABSVTX6 U77 ( .A(n61), .B(n954), .C(n953), .D(n952), .Z(n984) );
  AO6SVTX1 U78 ( .A(n1063), .B(m1[23]), .C(n1062), .Z(n1064) );
  IVSVTX2 U79 ( .A(n1548), .Z(n662) );
  NR2SVTX4 U80 ( .A(n978), .B(n977), .Z(n979) );
  AN2SVTX2 U81 ( .A(n65), .B(n847), .Z(n83) );
  AO6ABSVTX4 U82 ( .A(n648), .B(n647), .C(n71), .Z(n649) );
  ND4SVTX4 U83 ( .A(n1650), .B(n674), .C(n1113), .D(n794), .Z(n1321) );
  NR3SVTX2 U84 ( .A(n900), .B(n1664), .C(n882), .Z(n901) );
  AO7SVTX4 U85 ( .A(n912), .B(n913), .C(n911), .Z(n914) );
  ND2SVTX2 U86 ( .A(n1596), .B(n814), .Z(n815) );
  ND3ABSVTX2 U87 ( .A(n1053), .B(n1135), .C(n1051), .Z(n1055) );
  IVSVTX0H U88 ( .A(m1[24]), .Z(n1115) );
  AO3SVTX1 U89 ( .A(n957), .B(n1139), .C(n1061), .D(n1060), .Z(n502) );
  F_MUX21SVTX2 U90 ( .A(n24), .B(n25), .S(n1127), .Z(n648) );
  BFSVTX2 U91 ( .A(n963), .Z(n1051) );
  IVSVTX2 U92 ( .A(n609), .Z(n610) );
  ND3SVTX1 U93 ( .A(n725), .B(n724), .C(n795), .Z(n729) );
  F_MUX21NSVTX1 U94 ( .A(n829), .B(n828), .S(n827), .Z(n830) );
  IVSVTX0H U95 ( .A(n826), .Z(n823) );
  IVSVTX0H U96 ( .A(n925), .Z(n927) );
  IVSVTX0H U97 ( .A(n857), .Z(n860) );
  IVSVTX0H U98 ( .A(n846), .Z(n843) );
  AO7SVTX1 U99 ( .A(n853), .B(n852), .C(n851), .Z(n858) );
  NR2ASVTX4 U100 ( .A(n881), .B(n880), .Z(n885) );
  ND3SVTX2 U101 ( .A(n1092), .B(n518), .C(n519), .Z(n524) );
  MUX21NSVTX4 U102 ( .A(n910), .B(n909), .S(n908), .Z(n912) );
  ND4ABCSVTX4 U103 ( .A(n1075), .B(n1078), .C(n127), .D(n976), .Z(n978) );
  AO2ABSVTX4 U104 ( .C(n1296), .D(n402), .A(n779), .B(n1139), .Z(n403) );
  ND3SVTX1 U105 ( .A(n303), .B(n1239), .C(n1105), .Z(n1107) );
  IVSVTX2 U106 ( .A(n948), .Z(n937) );
  IVSVTX0H U107 ( .A(n693), .Z(n699) );
  IVSVTX0H U108 ( .A(n854), .Z(n856) );
  F_MUX21SVTX2 U109 ( .A(n645), .B(n644), .S(n26), .Z(n40) );
  ND3SVTX2 U110 ( .A(n1134), .B(n964), .C(n963), .Z(n970) );
  F_MUX21NSVTX1 U111 ( .A(n640), .B(n642), .S(n639), .Z(n646) );
  IVSVTX0H U112 ( .A(n787), .Z(n789) );
  IVSVTX0H U113 ( .A(n232), .Z(n742) );
  IVSVTX0H U114 ( .A(n866), .Z(n933) );
  ND2ASVTX4 U115 ( .A(n907), .B(n955), .Z(n908) );
  AO7SVTX1 U116 ( .A(n840), .B(n906), .C(n839), .Z(n845) );
  IVSVTX0H U117 ( .A(n869), .Z(n865) );
  IVSVTX4 U118 ( .A(n9), .Z(n873) );
  IVSVTX0H U119 ( .A(n844), .Z(n841) );
  AO7CSVTX2 U120 ( .A(n378), .B(n379), .C(n1139), .Z(n383) );
  NR2SVTX4 U121 ( .A(n594), .B(n593), .Z(n597) );
  AO7SVTX2 U122 ( .A(n895), .B(n894), .C(n893), .Z(n896) );
  ND3ABSVTX4 U123 ( .A(n52), .B(n53), .C(n579), .Z(n583) );
  AO7SVTX2 U124 ( .A(n520), .B(n861), .C(n1092), .Z(n521) );
  AO17SVTX1 U125 ( .A(n757), .B(n1620), .C(n756), .D(n755), .Z(n758) );
  NR2ASVTX2 U126 ( .A(n671), .B(n670), .Z(n773) );
  NR2ASVTX2 U127 ( .A(n497), .B(n496), .Z(n957) );
  IVSVTX6 U128 ( .A(n1094), .Z(n949) );
  IVSVTX2 U129 ( .A(n1127), .Z(n691) );
  IVSVTX6 U130 ( .A(n1491), .Z(n1238) );
  IVSVTX0H U131 ( .A(n882), .Z(n797) );
  IVSVTX0H U132 ( .A(n618), .Z(n619) );
  IVSVTX2 U133 ( .A(n1620), .Z(n1279) );
  IVSVTX2 U134 ( .A(n498), .Z(n958) );
  IVSVTX0H U135 ( .A(n695), .Z(n692) );
  CTIVSVTX2 U136 ( .A(n52), .Z(n10) );
  IVSVTX0H U137 ( .A(n849), .Z(n853) );
  IVSVTX0H U138 ( .A(n621), .Z(n810) );
  IVSVTX0H U139 ( .A(n965), .Z(n966) );
  IVSVTX0H U140 ( .A(n757), .Z(n754) );
  F_IVSVTX1 U141 ( .A(n57), .Z(n56) );
  IVSVTX0H U142 ( .A(n581), .Z(n53) );
  IVSVTX0H U143 ( .A(n881), .Z(n798) );
  CTIVSVTX8 U144 ( .A(n4), .Z(n1664) );
  CTIVSVTX8 U145 ( .A(n127), .Z(n4) );
  ND2SVTX2 U146 ( .A(m1[24]), .B(n534), .Z(n498) );
  IVSVTX8 U147 ( .A(n674), .Z(n1596) );
  IVSVTX0H U148 ( .A(n733), .Z(n685) );
  IVSVTX0H U149 ( .A(n690), .Z(n697) );
  IVSVTX0H U150 ( .A(n852), .Z(n782) );
  IVSVTX0H U151 ( .A(n836), .Z(n837) );
  IVSVTX0H U152 ( .A(n731), .Z(n732) );
  IVSVTX0H U153 ( .A(n676), .Z(n790) );
  IVSVTX0H U154 ( .A(n928), .Z(n864) );
  NR2ASVTX4 U155 ( .A(n819), .B(n826), .Z(n948) );
  IVSVTX0H U156 ( .A(n791), .Z(n677) );
  IVSVTX0H U157 ( .A(n1070), .Z(n400) );
  IVSVTX0H U158 ( .A(n548), .Z(n511) );
  ND2SVTX2 U159 ( .A(n543), .B(n542), .Z(n672) );
  BFSVTX8 U160 ( .A(n374), .Z(n1620) );
  IVSVTX0H U161 ( .A(n932), .Z(n930) );
  AO1SVTX2 U162 ( .A(n561), .B(n638), .C(n635), .D(n556), .Z(n559) );
  AO7NSVTX2 U163 ( .A(n545), .B(n512), .C(n546), .Z(n57) );
  IVSVTX2 U164 ( .A(n762), .Z(n315) );
  IVSVTX0H U165 ( .A(n745), .Z(n746) );
  IVSVTX0H U166 ( .A(n748), .Z(n751) );
  IVSVTX2 U167 ( .A(n568), .Z(n652) );
  IVSVTX0H U168 ( .A(n547), .Z(n512) );
  IVSVTX0H U169 ( .A(n735), .Z(n702) );
  IVSVTX0H U170 ( .A(n625), .Z(n626) );
  IVSVTX0H U171 ( .A(n749), .Z(n750) );
  F_IVSVTX1 U172 ( .A(n910), .Z(n905) );
  IVSVTX0H U173 ( .A(n1052), .Z(n362) );
  IVSVTX0H U174 ( .A(n1050), .Z(n363) );
  F_ND2ASVTX2 U175 ( .A(n359), .B(n1139), .Z(n1088) );
  CTAN2BSVTX4 U176 ( .A(n345), .B(n344), .Z(n1118) );
  AN2BSVTX2 U177 ( .A(n1138), .B(n305), .Z(n1087) );
  AO1CDSVTX4 U178 ( .A(n264), .B(n70), .C(n1109), .D(n1108), .Z(n261) );
  IVSVTX2 U179 ( .A(n636), .Z(n345) );
  NR2SVTX4 U180 ( .A(n852), .B(n555), .Z(n637) );
  AO7SVTX6 U181 ( .A(n259), .B(n531), .C(n258), .Z(n263) );
  ND3SVTX1 U182 ( .A(n539), .B(n1104), .C(n1105), .Z(n541) );
  OR2SVTX2 U183 ( .A(n889), .B(n895), .Z(n28) );
  OR2BSVTX4 U184 ( .A(n36), .B(m1[24]), .Z(n1108) );
  AO6SVTX4 U185 ( .A(n313), .B(n312), .C(n311), .Z(n1093) );
  ND2SVTX2 U186 ( .A(n447), .B(n446), .Z(n877) );
  B_ND2SVTX2 U187 ( .A(n463), .B(n675), .Z(n676) );
  IVSVTX2 U188 ( .A(n768), .Z(n771) );
  IVSVTX0H U189 ( .A(n538), .Z(n539) );
  IVSVTX2 U190 ( .A(n310), .Z(n93) );
  ND2SVTX4 U191 ( .A(n125), .B(n124), .Z(n312) );
  IVSVTX4 U192 ( .A(n429), .Z(n432) );
  B_ND2SVTX2 U193 ( .A(n748), .B(n372), .Z(n370) );
  OR2SVTX2 U194 ( .A(n1185), .B(n220), .Z(n330) );
  NR2SVTX2 U195 ( .A(m1[20]), .B(m1[23]), .Z(n618) );
  IVSVTX2 U196 ( .A(n32), .Z(n33) );
  AO6SVTX2 U197 ( .A(n395), .B(n63), .C(n394), .Z(n893) );
  NR2SVTX2 U198 ( .A(n359), .B(m1[22]), .Z(n965) );
  ND4SVTX1 U199 ( .A(m1[26]), .B(n1138), .C(m1[25]), .D(n1109), .Z(n326) );
  NR2ASVTX1 U200 ( .A(n117), .B(m1[22]), .Z(n255) );
  EOSVTX1 U201 ( .A(n1067), .B(n408), .Z(n453) );
  CTIVSVTX2 U202 ( .A(n398), .Z(n816) );
  NR2ASVTX2 U203 ( .A(n651), .B(m1[22]), .Z(n635) );
  ND2SVTX2 U204 ( .A(n359), .B(n535), .Z(n310) );
  IVSVTX0H U205 ( .A(n584), .Z(n585) );
  B_ND2SVTX2 U206 ( .A(n123), .B(n198), .Z(n124) );
  F_AN2SVTX2 U207 ( .A(n408), .B(n1136), .Z(n552) );
  AO6SVTX2 U208 ( .A(n1021), .B(n217), .C(n216), .Z(n218) );
  AN2SVTX4 U209 ( .A(n745), .B(n369), .Z(n372) );
  NR2SVTX2 U210 ( .A(n179), .B(n178), .Z(n1353) );
  ND2ASVTX6 U211 ( .A(n1635), .B(n1631), .Z(n177) );
  IVSVTX2 U212 ( .A(n230), .Z(n231) );
  F_AN2SVTX2 U213 ( .A(n296), .B(n117), .Z(n1359) );
  CTIVSVTX2 U214 ( .A(n337), .Z(n333) );
  B_ND2SVTX2 U215 ( .A(n462), .B(n342), .Z(n347) );
  OR2BSVTX4 U216 ( .A(n5), .B(m1[19]), .Z(n745) );
  AO7SVTX2 U217 ( .A(n1477), .B(n1474), .C(n1476), .Z(n1021) );
  B_ND2SVTX2 U218 ( .A(n140), .B(n1421), .Z(n995) );
  AN2SVTX4 U219 ( .A(n280), .B(n279), .Z(n281) );
  OR2SVTX2 U220 ( .A(m1[13]), .B(n277), .Z(n58) );
  EN3SVTX6 U221 ( .A(n1067), .B(m1[20]), .C(n534), .Z(n451) );
  ND2ASVTX4 U222 ( .A(m1[12]), .B(n433), .Z(n1652) );
  B_ND2SVTX2 U223 ( .A(n175), .B(n174), .Z(n1632) );
  ND2ASVTX6 U224 ( .A(n479), .B(n467), .Z(n8) );
  NR2ASVTX4 U225 ( .A(n173), .B(n172), .Z(n1635) );
  IVSVTX0H U226 ( .A(n35), .Z(n223) );
  FAS1SVTX2 U227 ( .A(m1[13]), .B(m1[16]), .CI(n433), .CO(n180), .Z(n178) );
  OR2BSVTX4 U228 ( .A(n31), .B(m1[14]), .Z(n1196) );
  NR2SVTX1 U229 ( .A(m1[23]), .B(n534), .Z(n203) );
  IVSVTX0H U230 ( .A(n283), .Z(n13) );
  ND2ASVTX4 U231 ( .A(m1[18]), .B(n463), .Z(n835) );
  F_ND2SVTX1 U232 ( .A(m1[19]), .B(n413), .Z(n349) );
  AO7SVTX2 U233 ( .A(n1495), .B(n1492), .C(n1494), .Z(n1003) );
  AO6SVTX2 U234 ( .A(n1513), .B(n1511), .C(n1510), .Z(n1575) );
  NR2SVTX2 U235 ( .A(m1[5]), .B(n276), .Z(n1474) );
  AO7SVTX2 U236 ( .A(n1647), .B(n1269), .C(n1270), .Z(n483) );
  AO7ABSVTX2 U237 ( .A(n1191), .B(n249), .C(n21), .Z(n20) );
  IVSVTX8 U238 ( .A(m1[23]), .Z(n1067) );
  IVSVTX0H U239 ( .A(n158), .Z(n138) );
  CTIVSVTX2 U240 ( .A(n174), .Z(n134) );
  IVSVTX0H U241 ( .A(n152), .Z(n142) );
  IVSVTX4 U242 ( .A(n169), .Z(n135) );
  ND2ASVTX4 U243 ( .A(m1[13]), .B(n433), .Z(n1284) );
  B_ND2SVTX2 U244 ( .A(m1[5]), .B(n285), .Z(n1494) );
  IVSVTX4 U245 ( .A(m1[27]), .Z(n1109) );
  IVSVTX0H U246 ( .A(n248), .Z(n233) );
  F_ND2ASVTX2 U247 ( .A(n293), .B(n296), .Z(n1176) );
  IVSVTX0H U248 ( .A(n1538), .Z(n145) );
  NR2SVTX2 U249 ( .A(m1[5]), .B(m1[2]), .Z(n1586) );
  AO7NSVTX1 U250 ( .A(n1615), .B(n67), .C(n1183), .Z(n21) );
  ND3ABSVTX4 U251 ( .A(m1[15]), .B(n96), .C(n408), .Z(n202) );
  B_ND2SVTX2 U252 ( .A(n277), .B(n276), .Z(n284) );
  CTIVSVTX10 U253 ( .A(n117), .Z(n5) );
  ND2ASVTX6 U254 ( .A(m1[17]), .B(n342), .Z(n253) );
  FAS1SVTX2 U255 ( .A(m1[5]), .B(n146), .CI(m1[6]), .CO(n155), .Z(n153) );
  IVSVTX0H U256 ( .A(n1467), .Z(n278) );
  FA1SVTX4 U257 ( .A(n7), .B(m1[12]), .CI(n31), .CO(n170), .Z(n167) );
  IVSVTX4 U258 ( .A(n532), .Z(n567) );
  ND4ABSVTX6 U259 ( .A(n87), .B(n96), .C(n97), .D(n16), .Z(n262) );
  IVSVTX2 U260 ( .A(m1[5]), .Z(n1487) );
  IVSVTX8 U261 ( .A(m1[21]), .Z(n532) );
  FAS1SVTX2 U262 ( .A(n285), .B(n31), .CI(n277), .CO(n168), .Z(n164) );
  IVSVTX2 U263 ( .A(m1[1]), .Z(n1523) );
  IVSVTX8 U264 ( .A(m1[17]), .Z(n413) );
  AN2SVTX4 U265 ( .A(n221), .B(n293), .Z(n16) );
  AN3SVTX4 U266 ( .A(n89), .B(n1371), .C(n117), .Z(n90) );
  IVSVTX8 U267 ( .A(n31), .Z(n293) );
  IVSVTX8 U268 ( .A(m1[16]), .Z(n117) );
  CTIVSVTX2 U269 ( .A(m1[6]), .Z(n103) );
  IVSVTX8 U270 ( .A(m1[15]), .Z(n316) );
  IVSVTX10 U271 ( .A(n89), .Z(n277) );
  IVSVTX4 U272 ( .A(n46), .Z(n47) );
  IVSVTX6 U273 ( .A(m1[8]), .Z(n1409) );
  IVSVTX6 U274 ( .A(m1[10]), .Z(n89) );
  IVSVTX4 U275 ( .A(m1[3]), .Z(n1572) );
  F_ND3SVTX2 U276 ( .A(n1409), .B(n103), .C(n187), .Z(n188) );
  F_IVSVTX0H U277 ( .A(n591), .Z(n592) );
  ND3ABSVTX1 U278 ( .A(n636), .B(n634), .C(n1119), .Z(n557) );
  IVSVTX0H U279 ( .A(n1087), .Z(n517) );
  F_ND2ASVTX2 U280 ( .A(m1[12]), .B(m1[14]), .Z(n1285) );
  ND2SVTX2 U281 ( .A(n534), .B(m1[23]), .Z(n229) );
  AO20SVTX4 U282 ( .A(n638), .B(n637), .C(n352), .D(n351), .Z(n1092) );
  IVSVTX0H U283 ( .A(n1481), .Z(n1483) );
  NR2SVTX0H U284 ( .A(n789), .B(n788), .Z(n793) );
  AO3SVTX1 U285 ( .A(n1092), .B(n1091), .C(n1090), .D(n1089), .Z(n1099) );
  NR2SVTX0H U286 ( .A(n1115), .B(n1114), .Z(n1116) );
  CTIVSVTX10 U287 ( .A(n1572), .Z(n146) );
  F_ND2SVTX0H U288 ( .A(n1615), .B(n1614), .Z(n1623) );
  AO17ASVTX2 U289 ( .A(n31), .B(n1274), .C(n1371), .D(n133), .Z(n175) );
  F_ND2SVTX0H U290 ( .A(n334), .B(n335), .Z(n228) );
  IVSVTX0H U291 ( .A(n884), .Z(n887) );
  F_ND2SVTX0H U292 ( .A(n1528), .B(n1527), .Z(n1529) );
  NR2SVTX2 U293 ( .A(m1[6]), .B(n1572), .Z(n1558) );
  F_ND2SVTX0H U294 ( .A(n1494), .B(n1493), .Z(n1500) );
  F_ND2SVTX0H U295 ( .A(n1426), .B(n1425), .Z(n1428) );
  NR2ASVTX1 U296 ( .A(n1387), .B(n1390), .Z(n998) );
  F_ND2SVTX0H U297 ( .A(n1209), .B(n1208), .Z(n1212) );
  ENSVTX0H U298 ( .A(n1194), .B(n1193), .Z(n1201) );
  IVSVTX0H U299 ( .A(n389), .Z(n119) );
  F_ND2SVTX0H U300 ( .A(n1632), .B(n1631), .Z(n1641) );
  IVSVTX4 U301 ( .A(n960), .Z(n974) );
  AO1SVTX1 U302 ( .A(n1296), .B(n1661), .C(n1660), .D(n1659), .Z(n1662) );
  AO6SVTX4 U303 ( .A(n1384), .B(n1381), .C(n1382), .Z(n1331) );
  F_ENSVTX2 U304 ( .A(n1322), .B(n1331), .Z(m2[17]) );
  IVSVTX2 U305 ( .A(n531), .Z(n1104) );
  IVSVTX2 U306 ( .A(n253), .Z(n683) );
  F_AN2SVTX2 U307 ( .A(n656), .B(n655), .Z(n1) );
  AN2SVTX4 U308 ( .A(n181), .B(n180), .Z(n2) );
  AN3SVTX4 U309 ( .A(n517), .B(n1085), .C(n353), .Z(n3) );
  AO7SVTX4 U310 ( .A(n718), .B(n717), .C(n716), .Z(n719) );
  IVSVTX2 U311 ( .A(n1150), .Z(n48) );
  ND2SVTX2 U312 ( .A(n1147), .B(n1146), .Z(n1148) );
  AO7SVTX2 U313 ( .A(n1664), .B(n1630), .C(n1629), .Z(m2[9]) );
  AO7SVTX2 U314 ( .A(n1238), .B(n1376), .C(n1375), .Z(n1377) );
  CTIVSVTX2 U315 ( .A(n1149), .Z(n1252) );
  ND3SVTX6 U316 ( .A(n403), .B(n405), .C(n404), .Z(n506) );
  ND2ASVTX4 U317 ( .A(n950), .B(n977), .Z(n951) );
  AO3CDSVTX1 U318 ( .A(n974), .B(n1601), .C(n1600), .D(n1599), .Z(m2[2]) );
  AO7SVTX2 U319 ( .A(n1238), .B(n1035), .C(n1034), .Z(n1036) );
  NR2ASVTX2 U320 ( .A(n4), .B(n794), .Z(n803) );
  AO7SVTX2 U321 ( .A(n1087), .B(n346), .C(n1088), .Z(n358) );
  NR3ABSVTX4 U322 ( .A(n971), .B(n970), .C(n969), .Z(n972) );
  IVSVTX2 U323 ( .A(n353), .Z(n346) );
  IVSVTX6 U324 ( .A(n566), .Z(n779) );
  AO7SVTX2 U325 ( .A(n1607), .B(n1606), .C(n1605), .Z(n1608) );
  CTIVSVTX2 U326 ( .A(n672), .Z(n673) );
  ND2SVTX8 U327 ( .A(n315), .B(n314), .Z(n566) );
  ND2SVTX4 U328 ( .A(n260), .B(n261), .Z(n527) );
  AO7SVTX2 U329 ( .A(n930), .B(n929), .C(n928), .Z(n931) );
  IVSVTX4 U330 ( .A(n22), .Z(n568) );
  IVSVTX4 U331 ( .A(n393), .Z(n1644) );
  F_ND2SVTX1 U332 ( .A(n6), .B(n548), .Z(n1070) );
  B_ND2SVTX2 U333 ( .A(n546), .B(n6), .Z(n550) );
  NR2SVTX2 U334 ( .A(n927), .B(n926), .Z(n935) );
  CTIVSVTX2 U335 ( .A(n1088), .Z(n1085) );
  IVSVTX4 U336 ( .A(n535), .Z(n540) );
  IVSVTX2 U337 ( .A(n447), .Z(n417) );
  ND2ASVTX4 U338 ( .A(n535), .B(n538), .Z(n768) );
  B_ND2SVTX2 U339 ( .A(n554), .B(n553), .Z(n558) );
  B_ND2SVTX2 U340 ( .A(n386), .B(n101), .Z(n122) );
  IVSVTX8 U341 ( .A(n651), .Z(n463) );
  B_ND2SVTX2 U342 ( .A(n1264), .B(n1263), .Z(n1268) );
  IVSVTX2 U343 ( .A(n453), .Z(n424) );
  NR2SVTX2 U344 ( .A(n68), .B(n1009), .Z(n1017) );
  CTIVSVTX2 U345 ( .A(n326), .Z(n329) );
  B_ND2SVTX1 U346 ( .A(n1394), .B(n1393), .Z(n1396) );
  B_ND2SVTX1 U347 ( .A(n1583), .B(n1582), .Z(n1588) );
  IVSVTX8 U348 ( .A(n1136), .Z(n1139) );
  IVSVTX10 U349 ( .A(n1409), .Z(n285) );
  NR2SVTX2 U350 ( .A(n1256), .B(n1255), .Z(n1257) );
  B_ND2SVTX2 U351 ( .A(n1167), .B(n1166), .Z(n1172) );
  B_ND2SVTX2 U352 ( .A(n1152), .B(n1151), .Z(n1153) );
  AO7SVTX2 U353 ( .A(n1664), .B(n1445), .C(n1444), .Z(m2[5]) );
  AO6ABSVTX4 U354 ( .A(n1319), .B(n1315), .C(n807), .Z(n808) );
  AO7SVTX2 U355 ( .A(n1664), .B(n1418), .C(n1417), .Z(m2[7]) );
  NR2SVTX2 U356 ( .A(n1302), .B(n1300), .Z(m2[26]) );
  NR2ASVTX4 U357 ( .A(n1252), .B(n1250), .Z(n1151) );
  ND2ASVTX6 U358 ( .A(n817), .B(n506), .Z(n1253) );
  AO7SVTX2 U359 ( .A(n1664), .B(n1663), .C(n1662), .Z(m2[11]) );
  IVSVTX4 U360 ( .A(n951), .Z(n952) );
  B_ND2SVTX2 U361 ( .A(n1258), .B(n1301), .Z(n1302) );
  CTIVSVTX2 U362 ( .A(n1258), .Z(n1299) );
  NR3SVTX4 U363 ( .A(n974), .B(n973), .C(n972), .Z(n980) );
  ND2SVTX4 U364 ( .A(n69), .B(n597), .Z(n598) );
  AO1CSVTX4 U365 ( .A(n72), .B(n1099), .C(n1098), .D(n1097), .Z(n1100) );
  ND2SVTX2 U366 ( .A(n678), .B(n873), .Z(n679) );
  ND3SVTX4 U367 ( .A(n1491), .B(n524), .C(n523), .Z(n954) );
  ND2ASVTX4 U368 ( .A(n1124), .B(n1132), .Z(n1300) );
  NR2ASVTX4 U369 ( .A(n567), .B(n779), .Z(n577) );
  F_ENSVTX2 U370 ( .A(n359), .B(n1117), .Z(n1123) );
  CTIVSVTX2 U371 ( .A(n379), .Z(n380) );
  IVSVTX2 U372 ( .A(n821), .Z(n801) );
  IVSVTX4 U373 ( .A(n573), .Z(n454) );
  CTIVSVTX2 U374 ( .A(n495), .Z(n496) );
  CTIVSVTX4 U375 ( .A(n372), .Z(n375) );
  AO6ASVTX6 U376 ( .A(n488), .B(n487), .C(n486), .Z(n489) );
  ND2ASVTX4 U377 ( .A(n555), .B(n343), .Z(n636) );
  IVSVTX2 U378 ( .A(n308), .Z(n95) );
  AO6SVTX2 U379 ( .A(n1481), .B(n1027), .C(n1026), .Z(n1435) );
  ND2ASVTX4 U380 ( .A(n450), .B(n23), .Z(n22) );
  AO6SVTX2 U381 ( .A(n483), .B(n470), .C(n482), .Z(n484) );
  IVSVTX4 U382 ( .A(n262), .Z(n301) );
  B_ND2SVTX1 U383 ( .A(n1643), .B(n1642), .Z(n1645) );
  IVSVTX4 U384 ( .A(n451), .Z(n23) );
  NR3SVTX2 U385 ( .A(n534), .B(n690), .C(n533), .Z(n537) );
  F_AN2SVTX2 U386 ( .A(n620), .B(n619), .Z(n84) );
  B_ND2SVTX2 U387 ( .A(n651), .B(n1139), .Z(n925) );
  FAS1SVTX2 U388 ( .A(n416), .B(n651), .CI(m1[19]), .CO(n447), .Z(n444) );
  B_ND2SVTX2 U389 ( .A(n651), .B(m1[22]), .Z(n625) );
  B_ND2SVTX1 U390 ( .A(n480), .B(n468), .Z(n252) );
  IVSVTX4 U391 ( .A(n20), .Z(n485) );
  AO7SVTX4 U392 ( .A(n1575), .B(n213), .C(n212), .Z(n214) );
  B_ND2SVTX1 U393 ( .A(n1402), .B(n1401), .Z(n1404) );
  F_ND2SVTX1 U394 ( .A(n1579), .B(n1578), .Z(n1593) );
  IVSVTX0H U395 ( .A(n811), .Z(n622) );
  CTIVSVTX2 U396 ( .A(n284), .Z(n1009) );
  B_ND2SVTX2 U397 ( .A(n398), .B(n117), .Z(n735) );
  IVSVTX0H U398 ( .A(n1028), .Z(n1029) );
  B_ND2SVTX2 U399 ( .A(n1476), .B(n1475), .Z(n1486) );
  B_ND2SVTX2 U400 ( .A(m1[19]), .B(m1[22]), .Z(n811) );
  F_IVSVTX1 U401 ( .A(n1393), .Z(n111) );
  IVSVTX8 U402 ( .A(n1067), .Z(n1136) );
  CTIVSVTX4 U403 ( .A(m1[19]), .Z(n398) );
  F_ND2SVTX1 U404 ( .A(n47), .B(m1[5]), .Z(n1579) );
  B_ND2SVTX2 U405 ( .A(n210), .B(n1573), .Z(n213) );
  CTIVSVTX2 U406 ( .A(n215), .Z(n209) );
  NR3ABSVTX4 U407 ( .A(n1155), .B(n1167), .C(n1159), .Z(n1156) );
  IVSVTX6 U408 ( .A(n1048), .Z(n41) );
  IVSVTX6 U409 ( .A(n1170), .Z(n1048) );
  AO7SVTX6 U410 ( .A(n1332), .B(n1331), .C(n1330), .Z(n1333) );
  AO2ASVTX6 U411 ( .C(n920), .D(n1312), .A(n1324), .B(n922), .Z(n923) );
  ND2SVTX6 U412 ( .A(n809), .B(n808), .Z(n924) );
  NR2ASVTX4 U413 ( .A(n1321), .B(n1320), .Z(n1382) );
  AO6SVTX2 U414 ( .A(n1596), .B(n1443), .C(n1442), .Z(n1444) );
  AO6SVTX2 U415 ( .A(n1296), .B(n1416), .C(n1415), .Z(n1417) );
  ENSVTX0H U416 ( .A(n1318), .B(n1307), .Z(m2[15]) );
  AO3SVTX1 U417 ( .A(n974), .B(n1509), .C(n1508), .D(n1507), .Z(m2[4]) );
  AO3SVTX1 U418 ( .A(n1664), .B(n1466), .C(n1465), .D(n1464), .Z(m2[3]) );
  AO3SVTX1 U419 ( .A(n1238), .B(n1536), .C(n1535), .D(n1534), .Z(m2[0]) );
  ND2SVTX4 U420 ( .A(n1306), .B(n1305), .Z(n1318) );
  ND3ABSVTX4 U421 ( .A(n887), .B(n1664), .C(n886), .Z(n1311) );
  AO1SVTX2 U422 ( .A(n1596), .B(n1235), .C(n1234), .D(n1233), .Z(n1236) );
  ND4SVTX6 U423 ( .A(n1103), .B(n1102), .C(n1101), .D(n1100), .Z(n1250) );
  AO3SVTX1 U424 ( .A(n1238), .B(n1557), .C(n1556), .D(n1555), .Z(m2[1]) );
  IVSVTX2 U425 ( .A(n1251), .Z(n1146) );
  ND2ASVTX4 U426 ( .A(n61), .B(n526), .Z(n986) );
  B_ND2SVTX1 U427 ( .A(n1039), .B(n1038), .Z(m2[6]) );
  AO7SVTX2 U428 ( .A(n503), .B(n502), .C(n501), .Z(n504) );
  ND3ABSVTX4 U429 ( .A(n1664), .B(n900), .C(n885), .Z(n1313) );
  ND3SVTX2 U430 ( .A(n1136), .B(n457), .C(n4), .Z(n458) );
  ND2ASVTX4 U431 ( .A(n680), .B(n679), .Z(n778) );
  AO6SVTX2 U432 ( .A(n1548), .B(n1037), .C(n1036), .Z(n1038) );
  ND3SVTX6 U433 ( .A(n876), .B(n875), .C(n874), .Z(n1324) );
  NR3ASVTX4 U434 ( .A(n613), .B(n1664), .C(n612), .Z(n614) );
  ND4ABCSVTX4 U435 ( .A(n944), .B(n127), .C(n661), .D(n660), .Z(n939) );
  NR2ASVTX6 U436 ( .A(n1596), .B(n551), .Z(n603) );
  F_ND2ASVTX2 U437 ( .A(n1080), .B(n654), .Z(n655) );
  NR3SVTX4 U438 ( .A(n1093), .B(n773), .C(n673), .Z(n794) );
  CTIVSVTX2 U439 ( .A(n37), .Z(n1095) );
  AO4SVTX4 U440 ( .A(n802), .B(n799), .C(n801), .D(n800), .Z(n1314) );
  AO6ABSVTX2 U441 ( .A(n1664), .B(n1008), .C(n85), .Z(n1039) );
  CTIVSVTX2 U442 ( .A(n975), .Z(n976) );
  ND2SVTX2 U443 ( .A(n381), .B(n380), .Z(n382) );
  IVSVTX10 U444 ( .A(n384), .Z(n1296) );
  AO6ASVTX4 U445 ( .A(n646), .B(n40), .C(n1238), .Z(n71) );
  B_ND2SVTX2 U446 ( .A(n1078), .B(n1075), .Z(n946) );
  IVSVTX10 U447 ( .A(n1596), .Z(n384) );
  NR2ASVTX4 U448 ( .A(n933), .B(n867), .Z(n870) );
  AO7ABSVTX6 U449 ( .A(n572), .B(n652), .C(n571), .Z(n609) );
  F_AN2SVTX2 U450 ( .A(n1596), .B(n1007), .Z(n85) );
  F_ENSVTX2 U451 ( .A(n813), .B(n812), .Z(n814) );
  F_IVSVTX1 U452 ( .A(n604), .Z(n605) );
  B_ND2SVTX2 U453 ( .A(n1113), .B(n1112), .Z(n1143) );
  B_ND2SVTX2 U454 ( .A(n1075), .B(n4), .Z(n950) );
  AO7SVTX4 U455 ( .A(n653), .B(n454), .C(n574), .Z(n1078) );
  CTIVSVTX2 U456 ( .A(n1238), .Z(n1122) );
  F_ENSVTX2 U457 ( .A(n761), .B(n760), .Z(n764) );
  F_IVSVTX1 U458 ( .A(n900), .Z(n883) );
  CTIVSVTX2 U459 ( .A(n828), .Z(n825) );
  ENSVTX0H U460 ( .A(n1032), .B(n1024), .Z(n1035) );
  IVSVTX4 U461 ( .A(n1093), .Z(n314) );
  B_ND2SVTX2 U462 ( .A(n562), .B(n560), .Z(n564) );
  NR2ASVTX2 U463 ( .A(n1139), .B(n378), .Z(n381) );
  AO7SVTX4 U464 ( .A(n33), .B(n1065), .C(n625), .Z(n591) );
  ND3SVTX1 U465 ( .A(n1139), .B(n498), .C(n495), .Z(n494) );
  B_ND2SVTX2 U466 ( .A(n653), .B(n652), .Z(n661) );
  CTIVSVTX2 U467 ( .A(n355), .Z(n354) );
  NR2ASVTX4 U468 ( .A(n516), .B(n1092), .Z(n355) );
  F_ND2SVTX1 U469 ( .A(n929), .B(n865), .Z(n868) );
  AO21DSVTX2 U470 ( .A(n1390), .B(n995), .C(n1503), .D(n1389), .Z(n1391) );
  IVSVTX10 U471 ( .A(n489), .Z(n955) );
  B_ND2SVTX2 U472 ( .A(n493), .B(n587), .Z(n495) );
  F_EOSVTX2 U473 ( .A(n1182), .B(n1181), .Z(n1204) );
  AO7SVTX2 U474 ( .A(n752), .B(n751), .C(n750), .Z(n756) );
  AO17SVTX2 U475 ( .A(n1104), .B(n537), .C(n536), .D(n535), .Z(n543) );
  IVSVTX2 U476 ( .A(n771), .Z(n49) );
  AO7SVTX6 U477 ( .A(n292), .B(n291), .C(n290), .Z(n374) );
  F_IVSVTX1 U478 ( .A(n352), .Z(n344) );
  NR3ABSVTX6 U479 ( .A(n1105), .B(n197), .C(n196), .Z(n208) );
  AO7SVTX6 U480 ( .A(n1634), .B(n177), .C(n176), .Z(n720) );
  IVSVTX2 U481 ( .A(n879), .Z(n418) );
  AO7SVTX6 U482 ( .A(n879), .B(n882), .C(n877), .Z(n827) );
  F_IVSVTX1 U483 ( .A(n877), .Z(n878) );
  ND2SVTX4 U484 ( .A(n93), .B(n666), .Z(n232) );
  AO6CSVTX4 U485 ( .A(n307), .B(n306), .C(m1[26]), .Z(n762) );
  CTIVSVTX2 U486 ( .A(n449), .Z(n410) );
  AO7SVTX6 U487 ( .A(n8), .B(n485), .C(n484), .Z(n486) );
  F_IVSVTX1 U488 ( .A(n835), .Z(n840) );
  F_IVSVTX1 U489 ( .A(n1063), .Z(n497) );
  IVSVTX2 U490 ( .A(n373), .Z(n744) );
  F_IVSVTX1 U491 ( .A(n558), .Z(n562) );
  CTIVSVTX2 U492 ( .A(n519), .Z(n522) );
  F_IVSVTX1 U493 ( .A(n711), .Z(n712) );
  NR2SVTX1 U494 ( .A(n545), .B(n511), .Z(n513) );
  B_ND2SVTX2 U495 ( .A(n961), .B(n964), .Z(n581) );
  AO6SVTX6 U496 ( .A(n1177), .B(n116), .C(n115), .Z(n393) );
  B_ND2SVTX2 U497 ( .A(n932), .B(n360), .Z(n365) );
  IVSVTX2 U498 ( .A(n444), .Z(n414) );
  BFSVTX2 U499 ( .A(n1020), .Z(n1478) );
  CTIVSVTX2 U500 ( .A(n1430), .Z(n1216) );
  B_ND2SVTX2 U501 ( .A(n967), .B(n966), .Z(n971) );
  ND2ASVTX6 U502 ( .A(n175), .B(n134), .Z(n1631) );
  NR2SVTX2 U503 ( .A(n1604), .B(n1603), .Z(n1609) );
  IVSVTX0H U504 ( .A(n1353), .Z(n1355) );
  NR2ASVTX4 U505 ( .A(n681), .B(n490), .Z(n906) );
  B_ND2SVTX2 U506 ( .A(n1348), .B(n1347), .Z(n1350) );
  AN2BSVTX4 U507 ( .A(n463), .B(n305), .Z(n634) );
  IVSVTX2 U508 ( .A(n995), .Z(n141) );
  F_IVSVTX1 U509 ( .A(n347), .Z(n855) );
  B_ND2SVTX2 U510 ( .A(n510), .B(n546), .Z(n399) );
  B_ND2SVTX2 U511 ( .A(n517), .B(n516), .Z(n519) );
  AO6SVTX2 U512 ( .A(n749), .B(n745), .C(n747), .Z(n371) );
  AO6SVTX6 U513 ( .A(n149), .B(n1542), .C(n1541), .Z(n1569) );
  AO6SVTX6 U514 ( .A(n733), .B(n349), .C(n348), .Z(n852) );
  NR2SVTX2 U515 ( .A(n1217), .B(n54), .Z(n280) );
  CTIVSVTX2 U516 ( .A(n681), .Z(n682) );
  B_ND2SVTX1 U517 ( .A(n736), .B(n735), .Z(n740) );
  CTIVSVTX2 U518 ( .A(n545), .Z(n6) );
  AO6SVTX4 U519 ( .A(n166), .B(n996), .C(n165), .Z(n430) );
  B_ND2SVTX2 U520 ( .A(m1[25]), .B(n534), .Z(n510) );
  IVSVTX0H U521 ( .A(n1643), .Z(n1266) );
  B_ND2SVTX1 U522 ( .A(n1568), .B(n1567), .Z(n1570) );
  B_ND2SVTX2 U523 ( .A(n179), .B(n178), .Z(n1352) );
  AO6SVTX6 U524 ( .A(n171), .B(n1602), .C(n1603), .Z(n1634) );
  IVSVTX4 U525 ( .A(n214), .Z(n1020) );
  AO7SVTX6 U526 ( .A(n109), .B(n1002), .C(n108), .Z(n1177) );
  NR3SVTX4 U527 ( .A(n1577), .B(n1591), .C(n1590), .Z(n473) );
  IVSVTX0H U528 ( .A(n1346), .Z(n1347) );
  F_IVSVTX1 U529 ( .A(n1084), .Z(n516) );
  AO6SVTX4 U530 ( .A(n105), .B(n1550), .C(n104), .Z(n1002) );
  IVSVTX0H U531 ( .A(n469), .Z(n1363) );
  CTIVSVTX2 U532 ( .A(n1176), .Z(n112) );
  AO7SVTX2 U533 ( .A(n1433), .B(n1018), .C(n1019), .Z(n216) );
  B_ND2SVTX2 U534 ( .A(m1[13]), .B(n5), .Z(n1264) );
  F_IVSVTX1 U535 ( .A(n326), .Z(n205) );
  B_ND2SVTX1 U536 ( .A(n1001), .B(n1000), .Z(n1006) );
  NR3ABSVTX4 U537 ( .A(n13), .B(n1274), .C(n191), .Z(n192) );
  CTIVSVTX2 U538 ( .A(n419), .Z(n420) );
  ND2ASVTX4 U539 ( .A(n173), .B(n172), .Z(n1633) );
  NR2ASVTX6 U540 ( .A(n170), .B(n135), .Z(n1603) );
  ND2ASVTX6 U541 ( .A(n170), .B(n135), .Z(n1602) );
  IVSVTX10 U542 ( .A(n88), .Z(n651) );
  IVSVTX10 U543 ( .A(n305), .Z(n534) );
  CTIVSVTX2 U544 ( .A(n1014), .Z(n279) );
  B_ND2SVTX1 U545 ( .A(n1495), .B(n1497), .Z(n1461) );
  B_ND2SVTX2 U546 ( .A(n1015), .B(n284), .Z(n1217) );
  IVSVTX2 U547 ( .A(n1210), .Z(n1394) );
  B_ND2SVTX1 U548 ( .A(n1610), .B(n58), .Z(n1612) );
  IVSVTX0H U549 ( .A(n1495), .Z(n1496) );
  ND2SVTX2 U550 ( .A(n242), .B(n1452), .Z(n1025) );
  IVSVTX0H U551 ( .A(n1424), .Z(n1425) );
  NR2SVTX2 U552 ( .A(n236), .B(n235), .Z(n237) );
  NR2SVTX1 U553 ( .A(n1429), .B(n282), .Z(n1431) );
  IVSVTX0H U554 ( .A(n1285), .Z(n1288) );
  IVSVTX0H U555 ( .A(n1286), .Z(n1287) );
  NR2SVTX4 U556 ( .A(n162), .B(n161), .Z(n1390) );
  IVSVTX4 U557 ( .A(m1[25]), .Z(n359) );
  IVSVTX8 U558 ( .A(m1[22]), .Z(n305) );
  IVSVTX2 U559 ( .A(n168), .Z(n136) );
  B_ND2SVTX1 U560 ( .A(n1584), .B(n1549), .Z(n1551) );
  F_IVSVTX1 U561 ( .A(n157), .Z(n139) );
  B_ND2SVTX2 U562 ( .A(m1[7]), .B(n38), .Z(n1019) );
  IVSVTX2 U563 ( .A(n132), .Z(n173) );
  ND2SVTX2 U564 ( .A(n1188), .B(n35), .Z(n220) );
  B_ND2SVTX2 U565 ( .A(n1619), .B(n1196), .Z(n1280) );
  AO6SVTX4 U566 ( .A(n1515), .B(n273), .C(n1514), .Z(n1563) );
  IVSVTX0H U567 ( .A(n1613), .Z(n1614) );
  IVSVTX0H U568 ( .A(n1561), .Z(n1562) );
  AO6SVTX2 U569 ( .A(n1561), .B(n1559), .C(n1558), .Z(n1010) );
  B_ND2SVTX2 U570 ( .A(n1559), .B(n1560), .Z(n1011) );
  IVSVTX2 U571 ( .A(n1517), .Z(n273) );
  B_ND2SVTX2 U572 ( .A(m1[2]), .B(n272), .Z(n1513) );
  IVSVTX4 U573 ( .A(m1[2]), .Z(n1545) );
  IVSVTX6 U574 ( .A(m1[4]), .Z(n1454) );
  IVSVTX12 U575 ( .A(n102), .Z(n7) );
  OR2SVTX4 U576 ( .A(n474), .B(n473), .Z(n1481) );
  AO7SVTX2 U577 ( .A(n474), .B(n473), .C(n472), .Z(n475) );
  CTIVSVTX4 U578 ( .A(n8), .Z(n478) );
  AO7SVTX2 U579 ( .A(n843), .B(n1127), .C(n842), .Z(n848) );
  IVSVTX8 U580 ( .A(n955), .Z(n1127) );
  ND2SVTX2 U581 ( .A(n31), .B(m1[13]), .Z(n1183) );
  IVSVTX2 U582 ( .A(n1341), .Z(n1342) );
  ND3SVTX2 U583 ( .A(n1248), .B(n1253), .C(n1341), .Z(n1249) );
  AO7SVTX4 U584 ( .A(n1162), .B(n1161), .C(n1327), .Z(n1046) );
  F_MUX21NSVTX1 U585 ( .A(n632), .B(n631), .S(n1065), .Z(n633) );
  ND2SVTX2 U586 ( .A(m1[19]), .B(n532), .Z(n854) );
  NR2SVTX2 U587 ( .A(n413), .B(m1[19]), .Z(n348) );
  AN2SVTX8 U588 ( .A(n527), .B(n578), .Z(n9) );
  IVSVTX10 U589 ( .A(n9), .Z(n960) );
  AN2SVTX4 U590 ( .A(n5), .B(n271), .Z(n733) );
  AO6ASVTX4 U591 ( .A(n365), .B(n871), .C(n361), .Z(n1140) );
  AO6ABSVTX6 U592 ( .A(n12), .B(n11), .C(n703), .Z(n704) );
  CTIVSVTX2 U593 ( .A(n1644), .Z(n11) );
  OR2SVTX4 U594 ( .A(n702), .B(n892), .Z(n12) );
  IVSVTX4 U595 ( .A(n1248), .Z(n1243) );
  IVSVTX8 U596 ( .A(m1[13]), .Z(n1274) );
  CTIVSVTX2 U597 ( .A(n1209), .Z(n110) );
  AO7ABSVTX4 U598 ( .A(m1[22]), .B(n566), .C(n947), .Z(n953) );
  ND4ASVTX8 U599 ( .A(n14), .B(n767), .C(n766), .D(n765), .Z(n1304) );
  AN2SVTX4 U600 ( .A(n65), .B(n734), .Z(n14) );
  OR2SVTX4 U601 ( .A(n316), .B(n416), .Z(n335) );
  NR3SVTX4 U602 ( .A(n282), .B(n1009), .C(n54), .Z(n289) );
  IVSVTX6 U603 ( .A(m1[9]), .Z(n102) );
  IVSVTX2 U604 ( .A(n527), .Z(n818) );
  ND3SVTX4 U605 ( .A(n873), .B(n79), .C(n872), .Z(n874) );
  OR2SVTX4 U606 ( .A(n868), .B(n870), .Z(n79) );
  ND3SVTX6 U607 ( .A(n198), .B(n123), .C(n301), .Z(n230) );
  IVSVTX4 U608 ( .A(n198), .Z(n200) );
  AO6SVTX2 U609 ( .A(n1397), .B(n1214), .C(n1213), .Z(n286) );
  AO7SVTX6 U610 ( .A(n1569), .B(n428), .C(n427), .Z(n429) );
  AO6CSVTX4 U611 ( .A(n66), .B(n400), .C(n1114), .Z(n401) );
  IVSVTX8 U612 ( .A(n27), .Z(n66) );
  F_ND2ASVTX2 U613 ( .A(n316), .B(n271), .Z(n366) );
  AN2SVTX2 U614 ( .A(n355), .B(n1088), .Z(n15) );
  NR2SVTX2 U615 ( .A(n15), .B(n1238), .Z(n356) );
  AO7SVTX8 U616 ( .A(n219), .B(n1020), .C(n218), .Z(n1403) );
  F_AN2SVTX2 U617 ( .A(n146), .B(n1487), .Z(n75) );
  IVSVTX4 U618 ( .A(n1140), .Z(n52) );
  CTIVSVTX2 U619 ( .A(n969), .Z(n968) );
  AO7SVTX2 U620 ( .A(n676), .B(n788), .C(n787), .Z(n871) );
  IVSVTX6 U621 ( .A(m1[12]), .Z(n221) );
  AO1SVTX4 U622 ( .A(n698), .B(n1127), .C(n17), .D(n232), .Z(n19) );
  AO2NSVTX2 U623 ( .A(n698), .B(n697), .C(n696), .D(n695), .Z(n17) );
  NR2ASVTX4 U624 ( .A(n694), .B(n695), .Z(n698) );
  F_IVSVTX0H U625 ( .A(n769), .Z(n770) );
  ND4ASVTX4 U626 ( .A(n36), .B(n304), .C(n1138), .D(n266), .Z(n267) );
  NR2SVTX2 U627 ( .A(n163), .B(n164), .Z(n18) );
  F_EOSVTX2 U628 ( .A(n1139), .B(n401), .Z(n402) );
  NR2SVTX0H U629 ( .A(n1067), .B(n1070), .Z(n1073) );
  AO6SVTX4 U630 ( .A(n289), .B(n1012), .C(n288), .Z(n290) );
  F_AN2SVTX2 U631 ( .A(n89), .B(m1[7]), .Z(n68) );
  AO7SVTX2 U632 ( .A(n1406), .B(n248), .C(n247), .Z(n1191) );
  IVSVTX2 U633 ( .A(n1106), .Z(n195) );
  NR3SVTX2 U634 ( .A(n531), .B(n1107), .C(n1106), .Z(n1111) );
  ND2SVTX2 U635 ( .A(n1602), .B(n137), .Z(n1173) );
  IVSVTX2 U636 ( .A(n1607), .Z(n137) );
  CTIVSVTX2 U637 ( .A(n468), .Z(n481) );
  AO7SVTX4 U638 ( .A(n287), .B(n1215), .C(n286), .Z(n288) );
  AN3SVTX4 U639 ( .A(n1313), .B(n1312), .C(n1311), .Z(n1332) );
  IVSVTX2 U640 ( .A(n331), .Z(n332) );
  ND2SVTX2 U641 ( .A(n1284), .B(n1285), .Z(n331) );
  IVSVTX4 U642 ( .A(n850), .Z(n343) );
  NR2SVTX2 U643 ( .A(n850), .B(n853), .Z(n857) );
  AO6ABSVTX4 U644 ( .A(n1401), .B(n55), .C(n1221), .Z(n1184) );
  AO6SVTX4 U645 ( .A(n781), .B(n780), .C(n81), .Z(n785) );
  ND2SVTX4 U646 ( .A(n276), .B(n1030), .Z(n96) );
  CTIVSVTX2 U647 ( .A(n1030), .Z(n239) );
  CTIVSVTX2 U648 ( .A(n1222), .Z(n55) );
  ND2SVTX2 U649 ( .A(n31), .B(n102), .Z(n1222) );
  AO7SVTX4 U650 ( .A(n114), .B(n1178), .C(n113), .Z(n115) );
  AO6SVTX4 U651 ( .A(n64), .B(n1180), .C(n112), .Z(n113) );
  IVSVTX2 U652 ( .A(n1610), .Z(n1180) );
  AO17SVTX2 U653 ( .A(n459), .B(n1094), .C(n458), .D(n817), .Z(n1254) );
  ND3SVTX2 U654 ( .A(n611), .B(n605), .C(n1094), .Z(n608) );
  ND3SVTX2 U655 ( .A(n1121), .B(n760), .C(n1118), .Z(n1090) );
  ND3SVTX4 U656 ( .A(n689), .B(n1491), .C(n688), .Z(n708) );
  CTIVSVTX2 U657 ( .A(n492), .Z(n465) );
  CTIVSVTX2 U658 ( .A(n1125), .Z(n1126) );
  ND3SVTX4 U659 ( .A(n558), .B(n559), .C(n557), .Z(n565) );
  AO3SVTX6 U660 ( .A(n295), .B(n1278), .C(n294), .D(n1276), .Z(n748) );
  ND2SVTX2 U661 ( .A(m1[15]), .B(m1[13]), .Z(n1270) );
  IVSVTX4 U662 ( .A(n752), .Z(n369) );
  OR2SVTX8 U663 ( .A(m1[15]), .B(n271), .Z(n368) );
  IVSVTX6 U664 ( .A(n915), .Z(n1308) );
  ND3ABSVTX6 U665 ( .A(n818), .B(n1093), .C(n1308), .Z(n606) );
  NR2SVTX2 U666 ( .A(n838), .B(n837), .Z(n844) );
  IVSVTX10 U667 ( .A(n532), .Z(n462) );
  B_ND2SVTX2 U668 ( .A(n958), .B(n956), .Z(n959) );
  F_ND3SVTX2 U669 ( .A(n918), .B(n917), .C(n1310), .Z(n919) );
  ND2SVTX4 U670 ( .A(n333), .B(n332), .Z(n340) );
  OR2SVTX2 U671 ( .A(n398), .B(m1[22]), .Z(n928) );
  IVSVTX4 U672 ( .A(n606), .Z(n607) );
  IVSVTX4 U673 ( .A(n177), .Z(n710) );
  ND2SVTX4 U674 ( .A(n1320), .B(n1319), .Z(n1381) );
  AO7SVTX2 U675 ( .A(n250), .B(n1407), .C(n485), .Z(n1648) );
  AO6CSVTX4 U676 ( .A(n963), .B(n791), .C(n676), .Z(n792) );
  IVSVTX2 U677 ( .A(n962), .Z(n964) );
  NR2SVTX2 U678 ( .A(m1[8]), .B(m1[6]), .Z(n1030) );
  ND2SVTX2 U679 ( .A(n1405), .B(n233), .Z(n1192) );
  ENSVTX4 U680 ( .A(n1339), .B(n1338), .Z(m2[19]) );
  CTIVSVTX2 U681 ( .A(n632), .Z(n628) );
  AO7SVTX2 U682 ( .A(n1664), .B(n1206), .C(n1205), .Z(m2[10]) );
  AO6ABSVTX2 U683 ( .A(n1192), .B(n1407), .C(n1191), .Z(n1616) );
  IVSVTX4 U684 ( .A(m1[7]), .Z(n276) );
  AO7SVTX4 U685 ( .A(n1303), .B(n1304), .C(n1317), .Z(n774) );
  ND3SVTX2 U686 ( .A(n873), .B(n1059), .C(n1058), .Z(n1103) );
  ND3SVTX2 U687 ( .A(m1[24]), .B(n1055), .C(n1054), .Z(n1059) );
  AO6SVTX4 U688 ( .A(n107), .B(n1003), .C(n106), .Z(n108) );
  IVSVTX4 U689 ( .A(n834), .Z(n922) );
  ND2SVTX4 U690 ( .A(n445), .B(n444), .Z(n882) );
  FAS1SVTX4 U691 ( .A(m1[7]), .B(n277), .CI(n7), .CO(n163), .Z(n162) );
  AO7SVTX4 U692 ( .A(n1258), .B(n1249), .C(n1300), .Z(n43) );
  ND2SVTX4 U693 ( .A(n527), .B(n578), .Z(n1548) );
  AO6SVTX4 U694 ( .A(n66), .B(n513), .C(n56), .Z(n514) );
  ND2SVTX2 U695 ( .A(m1[20]), .B(m1[23]), .Z(n620) );
  IVSVTX2 U696 ( .A(n1010), .Z(n275) );
  NR2SVTX2 U697 ( .A(n687), .B(n686), .Z(n688) );
  ND2SVTX2 U698 ( .A(n1359), .B(n334), .Z(n336) );
  NR3SVTX6 U699 ( .A(n1259), .B(n43), .C(n44), .Z(m2[25]) );
  NR2ASVTX2 U700 ( .A(n1136), .B(n1075), .Z(n1077) );
  OR2SVTX4 U701 ( .A(n293), .B(n1274), .Z(n133) );
  AO5ASVTX2 U702 ( .B(n408), .A(m1[19]), .C(n305), .Z(n450) );
  ND2SVTX2 U703 ( .A(n1160), .B(n1040), .Z(n1341) );
  F_ND3SVTX2 U704 ( .A(n960), .B(n916), .C(n915), .Z(n805) );
  ND2SVTX2 U705 ( .A(n327), .B(n205), .Z(n206) );
  AO7SVTX2 U706 ( .A(n1426), .B(n999), .C(n1001), .Z(n106) );
  BFSVTX12 U707 ( .A(m1[11]), .Z(n31) );
  F_ND2ASVTX2 U708 ( .A(m1[7]), .B(n1487), .Z(n242) );
  AO7ABSVTX6 U709 ( .A(n1248), .B(n1044), .C(n1043), .Z(n1170) );
  IVSVTX8 U710 ( .A(m1[20]), .Z(n88) );
  NR2SVTX2 U711 ( .A(n1085), .B(n1084), .Z(n1121) );
  NR2SVTX2 U712 ( .A(n938), .B(n937), .Z(n940) );
  ND2SVTX2 U713 ( .A(n4), .B(n661), .Z(n938) );
  ND2SVTX2 U714 ( .A(n1049), .B(n974), .Z(n1149) );
  NR2SVTX2 U715 ( .A(n864), .B(n930), .Z(n869) );
  F_ND2ASVTX2 U716 ( .A(m1[19]), .B(m1[22]), .Z(n932) );
  ND2SVTX2 U717 ( .A(n1052), .B(n1136), .Z(n1137) );
  ND2SVTX4 U718 ( .A(n1327), .B(n1247), .Z(n1339) );
  AO7SVTX2 U719 ( .A(n871), .B(n870), .C(n869), .Z(n872) );
  AO7NSVTX2 U720 ( .A(n1086), .B(n1090), .C(n1491), .Z(n72) );
  AN2BSVTX4 U721 ( .A(n209), .B(n283), .Z(n1479) );
  IVSVTX10 U722 ( .A(m1[24]), .Z(n1138) );
  FAS1SVTX4 U723 ( .A(m1[22]), .B(m1[24]), .CI(m1[25]), .Z(n419) );
  ND2SVTX2 U724 ( .A(n462), .B(m1[24]), .Z(n546) );
  ND3ABSVTX4 U725 ( .A(n697), .B(n692), .C(n691), .Z(n700) );
  ND2SVTX2 U726 ( .A(n239), .B(n241), .Z(n245) );
  IVSVTX2 U727 ( .A(n238), .Z(n241) );
  ND2SVTX2 U728 ( .A(n296), .B(n413), .Z(n1367) );
  ND3SVTX4 U729 ( .A(n760), .B(n1118), .C(n516), .Z(n353) );
  ND2SVTX4 U730 ( .A(n508), .B(n507), .Z(n509) );
  ND2SVTX2 U731 ( .A(n534), .B(n422), .Z(n423) );
  ND2SVTX4 U732 ( .A(n451), .B(n450), .Z(n653) );
  IVSVTX2 U733 ( .A(n364), .Z(n788) );
  IVSVTX2 U734 ( .A(n871), .Z(n929) );
  ND2SVTX2 U735 ( .A(n567), .B(n271), .Z(n364) );
  ND3SVTX4 U736 ( .A(n700), .B(n699), .C(n19), .Z(n707) );
  F_ENSVTX2 U737 ( .A(n82), .B(n704), .Z(n705) );
  ND2SVTX2 U738 ( .A(m1[13]), .B(n277), .Z(n1610) );
  NR2ASVTX2 U739 ( .A(n272), .B(n1572), .Z(n1517) );
  IVSVTX4 U740 ( .A(m1[0]), .Z(n272) );
  ND3SVTX4 U741 ( .A(n544), .B(n672), .C(n578), .Z(n915) );
  B_ND2SVTX1 U742 ( .A(n828), .B(n826), .Z(n829) );
  ND2SVTX2 U743 ( .A(n820), .B(n819), .Z(n828) );
  AO7SVTX4 U744 ( .A(n456), .B(n1080), .C(n455), .Z(n499) );
  ND2SVTX2 U745 ( .A(n296), .B(m1[16]), .Z(n1364) );
  ND2SVTX4 U746 ( .A(n334), .B(n1360), .Z(n337) );
  AO3SVTX2 U747 ( .A(n338), .B(n337), .C(n336), .D(n335), .Z(n339) );
  IVSVTX4 U748 ( .A(n957), .Z(n1130) );
  ND2SVTX2 U749 ( .A(m1[19]), .B(n567), .Z(n836) );
  AO6SVTX6 U750 ( .A(n1343), .B(n1342), .C(n985), .Z(n1344) );
  ND2SVTX2 U751 ( .A(m1[18]), .B(n463), .Z(n851) );
  NR2SVTX2 U752 ( .A(n638), .B(n637), .Z(n641) );
  AO7SVTX2 U753 ( .A(n1053), .B(n1140), .C(n1137), .Z(n1057) );
  IVSVTX4 U754 ( .A(n1321), .Z(n1319) );
  AN2SVTX4 U755 ( .A(n574), .B(n573), .Z(n78) );
  ND2SVTX2 U756 ( .A(n453), .B(n452), .Z(n574) );
  ND2ASVTX8 U757 ( .A(n452), .B(n424), .Z(n573) );
  AO7ABSVTX2 U758 ( .A(m1[23]), .B(m1[20]), .C(n423), .Z(n452) );
  NR2SVTX2 U759 ( .A(n1538), .B(n237), .Z(n1590) );
  NR2SVTX2 U760 ( .A(m1[5]), .B(n47), .Z(n1577) );
  IVSVTX2 U761 ( .A(n282), .Z(n1015) );
  NR2SVTX2 U762 ( .A(n102), .B(m1[6]), .Z(n282) );
  AO7SVTX4 U763 ( .A(n906), .B(n492), .C(n491), .Z(n587) );
  B_ND2SVTX1 U764 ( .A(n906), .B(n910), .Z(n909) );
  IVSVTX0H U765 ( .A(n906), .Z(n904) );
  ND2SVTX2 U766 ( .A(m1[23]), .B(n1050), .Z(n1053) );
  NR2SVTX2 U767 ( .A(n962), .B(n965), .Z(n1050) );
  AO7SVTX2 U768 ( .A(n1664), .B(n1316), .C(n1315), .Z(n1384) );
  ND2SVTX4 U769 ( .A(n1318), .B(n1317), .Z(n1320) );
  ND2SVTX2 U770 ( .A(n1277), .B(n1651), .Z(n294) );
  ND2SVTX4 U771 ( .A(n795), .B(n796), .Z(n657) );
  AO6ABSVTX2 U772 ( .A(n211), .B(n1574), .C(n75), .Z(n212) );
  AO6SVTX2 U773 ( .A(n284), .B(n1429), .C(n68), .Z(n1215) );
  IVSVTX4 U774 ( .A(n341), .Z(n226) );
  AO7ABSVTX4 U775 ( .A(n1633), .B(n1632), .C(n1631), .Z(n176) );
  AO7SVTX4 U776 ( .A(n889), .B(n893), .C(n891), .Z(n396) );
  AO6SVTX1 U777 ( .A(n1498), .B(n1004), .C(n1003), .Z(n1427) );
  IVSVTX4 U778 ( .A(n390), .Z(n392) );
  AO7SVTX2 U779 ( .A(n702), .B(n894), .C(n736), .Z(n703) );
  IVSVTX4 U780 ( .A(n737), .Z(n894) );
  NR2SVTX2 U781 ( .A(n1479), .B(n1474), .Z(n1022) );
  NR2SVTX2 U782 ( .A(n295), .B(n1280), .Z(n373) );
  CTIVSVTX2 U783 ( .A(n819), .Z(n569) );
  AO6SVTX2 U784 ( .A(n66), .B(n810), .C(n622), .Z(n623) );
  ND3ABSVTX4 U785 ( .A(n33), .B(n629), .C(n955), .Z(n595) );
  CTIVSVTX2 U786 ( .A(n552), .Z(n554) );
  AN2SVTX0H U787 ( .A(n7), .B(m1[7]), .Z(n240) );
  NR2SVTX2 U788 ( .A(n1664), .B(n1136), .Z(n500) );
  AO6SVTX2 U789 ( .A(n1648), .B(n467), .C(n483), .Z(n1365) );
  CTIVSVTX2 U790 ( .A(n726), .Z(n724) );
  IVSVTX6 U791 ( .A(n65), .Z(n1650) );
  CTIVSVTX2 U792 ( .A(n635), .Z(n350) );
  IVSVTX2 U793 ( .A(n1223), .Z(n1401) );
  EO3SVTX4 U794 ( .A(m1[13]), .B(n31), .C(n296), .Z(n172) );
  CTIVSVTX4 U795 ( .A(n1173), .Z(n1639) );
  IVSVTX4 U796 ( .A(n1605), .Z(n171) );
  F_ND2ASVTX1 U797 ( .A(n1519), .B(n1518), .Z(n1520) );
  ENSVTX0H U798 ( .A(n1517), .B(n1516), .Z(n1525) );
  F_ND2SVTX0H U799 ( .A(n1176), .B(n64), .Z(n1182) );
  AO4SVTX1 U800 ( .A(n974), .B(n317), .C(n39), .D(n316), .Z(n318) );
  ND2SVTX2 U801 ( .A(n1251), .B(n1250), .Z(n1256) );
  AO1CDSVTX2 U802 ( .A(n1254), .B(n988), .C(n1253), .D(n1252), .Z(n1255) );
  ND2SVTX2 U803 ( .A(n1398), .B(n1214), .Z(n54) );
  AO7SVTX1 U804 ( .A(n433), .B(m1[18]), .C(n416), .Z(n434) );
  IVSVTX0H U805 ( .A(n642), .Z(n643) );
  CTIVSVTX2 U806 ( .A(n641), .Z(n639) );
  F_ND2SVTX0H U807 ( .A(n636), .B(n642), .Z(n640) );
  B_ND2SVTX1 U808 ( .A(n641), .B(n642), .Z(n645) );
  AO7SVTX2 U809 ( .A(n1364), .B(n481), .C(n480), .Z(n482) );
  IVSVTX0H U810 ( .A(n694), .Z(n696) );
  ND4ABSVTX2 U811 ( .A(n651), .B(n462), .C(n683), .D(n1139), .Z(n533) );
  ND2SVTX2 U812 ( .A(m1[18]), .B(n651), .Z(n839) );
  AO7SVTX2 U813 ( .A(n363), .B(n1140), .C(n362), .Z(n378) );
  F_ND2ASVTX2 U814 ( .A(n651), .B(m1[23]), .Z(n360) );
  AO7SVTX2 U815 ( .A(n367), .B(n1367), .C(n366), .Z(n749) );
  CTIVSVTX2 U816 ( .A(n210), .Z(n211) );
  NR2SVTX2 U817 ( .A(n1563), .B(n1011), .Z(n274) );
  F_ND2SVTX0H U818 ( .A(n31), .B(n1274), .Z(n222) );
  IVSVTX2 U819 ( .A(n717), .Z(n715) );
  AN2SVTX4 U820 ( .A(n304), .B(n303), .Z(n300) );
  NR2SVTX2 U821 ( .A(n910), .B(n343), .Z(n783) );
  IVSVTX2 U822 ( .A(n938), .Z(n654) );
  AO7SVTX2 U823 ( .A(n811), .B(n618), .C(n620), .Z(n547) );
  NR2SVTX2 U824 ( .A(n462), .B(m1[24]), .Z(n545) );
  ND2SVTX2 U825 ( .A(n466), .B(n465), .Z(n629) );
  IVSVTX2 U826 ( .A(n448), .Z(n409) );
  NR2SVTX2 U827 ( .A(n1138), .B(n567), .Z(n962) );
  B_ND2SVTX0H U828 ( .A(n462), .B(m1[23]), .Z(n421) );
  F_IVSVTX0H U829 ( .A(n1061), .Z(n1062) );
  F_ND2SVTX0H U830 ( .A(m1[18]), .B(n532), .Z(n787) );
  OR2SVTX0H U831 ( .A(n790), .B(n677), .Z(n62) );
  ND2SVTX2 U832 ( .A(n684), .B(n26), .Z(n689) );
  NR2SVTX0H U833 ( .A(n840), .B(n907), .Z(n846) );
  IVSVTX2 U834 ( .A(n760), .Z(n861) );
  NR2SVTX0H U835 ( .A(n856), .B(n855), .Z(n859) );
  IVSVTX2 U836 ( .A(n963), .Z(n867) );
  IVSVTX2 U837 ( .A(n360), .Z(n926) );
  AO7SVTX1 U838 ( .A(n961), .B(n965), .C(n967), .Z(n1052) );
  AO7SVTX2 U839 ( .A(n1530), .B(n1526), .C(n1528), .Z(n1550) );
  CTIVSVTX4 U840 ( .A(m1[3]), .Z(n46) );
  NR2SVTX2 U841 ( .A(m1[6]), .B(n146), .Z(n1581) );
  ND2SVTX4 U842 ( .A(n1067), .B(n463), .Z(n422) );
  AO7SVTX2 U843 ( .A(n1589), .B(n1577), .C(n1579), .Z(n474) );
  F_ND2ASVTX1 U844 ( .A(m1[6]), .B(n1454), .Z(n1452) );
  F_ND2SVTX0H U845 ( .A(m1[7]), .B(n1454), .Z(n1458) );
  AN2SVTX0H U846 ( .A(n285), .B(m1[6]), .Z(n1028) );
  IVSVTX2 U847 ( .A(m1[6]), .Z(n215) );
  NR2SVTX2 U848 ( .A(n1390), .B(n1385), .Z(n166) );
  AN2SVTX4 U849 ( .A(n1274), .B(n293), .Z(n67) );
  AO6SVTX2 U850 ( .A(n1286), .B(n1284), .C(n1283), .Z(n338) );
  ND2SVTX2 U851 ( .A(n675), .B(n316), .Z(n334) );
  ND2SVTX2 U852 ( .A(n129), .B(n128), .Z(n131) );
  F_ND2SVTX0H U853 ( .A(n296), .B(n675), .Z(n129) );
  NR2SVTX2 U854 ( .A(n1067), .B(n1239), .Z(n258) );
  F_ENSVTX2 U855 ( .A(n761), .B(n955), .Z(n734) );
  F_EOSVTX2 U856 ( .A(n740), .B(n739), .Z(n741) );
  AO6SVTX2 U857 ( .A(n95), .B(n94), .C(n93), .Z(n743) );
  F_ND2ASVTX2 U858 ( .A(n78), .B(n4), .Z(n604) );
  AO8SVTX2 U859 ( .A(n933), .B(n932), .C(n963), .D(n931), .Z(n934) );
  ND2SVTX2 U860 ( .A(n1296), .B(n624), .Z(n650) );
  AO6SVTX2 U861 ( .A(n66), .B(n548), .C(n547), .Z(n549) );
  IVSVTX2 U862 ( .A(n943), .Z(n1075) );
  F_ND2ASVTX2 U863 ( .A(m1[25]), .B(n534), .Z(n967) );
  AO7SVTX2 U864 ( .A(n962), .B(n1140), .C(n961), .Z(n969) );
  NR2SVTX2 U865 ( .A(n461), .B(n460), .Z(n505) );
  F_ND2ASVTX2 U866 ( .A(n1139), .B(n958), .Z(n1061) );
  AO6SVTX1 U867 ( .A(n1088), .B(n1087), .C(n1120), .Z(n1089) );
  B_ND2SVTX0H U868 ( .A(m1[24]), .B(n1093), .Z(n1098) );
  IVSVTX2 U869 ( .A(n1055), .Z(n1056) );
  F_ENSVTX2 U870 ( .A(n793), .B(n792), .Z(n916) );
  F_ND2SVTX0H U871 ( .A(n891), .B(n890), .Z(n899) );
  IVSVTX0H U872 ( .A(n889), .Z(n890) );
  NR2SVTX2 U873 ( .A(n530), .B(n529), .Z(n544) );
  NR2SVTX2 U874 ( .A(n1239), .B(n769), .Z(n530) );
  NR2ASVTX1 U875 ( .A(n841), .B(n845), .Z(n842) );
  AO3CDSVTX1 U876 ( .A(n861), .B(n860), .C(n859), .D(n858), .Z(n862) );
  ND2SVTX2 U877 ( .A(n194), .B(n408), .Z(n1106) );
  IVSVTX2 U878 ( .A(n1134), .Z(n1135) );
  NR2SVTX2 U879 ( .A(n1531), .B(n283), .Z(n1519) );
  F_AN2SVTX2 U880 ( .A(m1[1]), .B(n47), .Z(n1538) );
  IVSVTX0H U881 ( .A(n1581), .Z(n1582) );
  F_ND2ASVTX2 U882 ( .A(n1454), .B(n1545), .Z(n1573) );
  IVSVTX2 U883 ( .A(n153), .Z(n143) );
  FAS1SVTX2 U884 ( .A(m1[7]), .B(n285), .CI(m1[5]), .CO(n159), .Z(n157) );
  AO7SVTX1 U885 ( .A(n1030), .B(n1435), .C(n1029), .Z(n1031) );
  AO7SVTX2 U886 ( .A(n1014), .B(n1470), .C(n1013), .Z(n1430) );
  F_ND2SVTX0H U887 ( .A(n1406), .B(n1405), .Z(n1408) );
  AO7SVTX1 U888 ( .A(n1613), .B(n1616), .C(n1615), .Z(n1193) );
  OR2SVTX2 U889 ( .A(n31), .B(n296), .Z(n64) );
  F_ND2SVTX0H U890 ( .A(n1277), .B(n1276), .Z(n1282) );
  ND2SVTX2 U891 ( .A(n5), .B(n1371), .Z(n1360) );
  F_ND2SVTX0H U892 ( .A(n1368), .B(n1367), .Z(n1370) );
  F_ND2ASVTX2 U893 ( .A(n1265), .B(n1263), .Z(n391) );
  ENSVTX0H U894 ( .A(n299), .B(n298), .Z(n317) );
  NR2ASVTX1 U895 ( .A(n366), .B(n367), .Z(n299) );
  IVSVTX0H U896 ( .A(n1368), .Z(n297) );
  ND2SVTX2 U897 ( .A(n131), .B(n130), .Z(n716) );
  IVSVTX2 U898 ( .A(n66), .Z(n812) );
  AN3SVTX2 U899 ( .A(n78), .B(n653), .C(n610), .Z(n613) );
  MUX21NSVTX2 U900 ( .A(n959), .B(n958), .S(n1130), .Z(n981) );
  NR2SVTX2 U901 ( .A(n778), .B(n777), .Z(n1315) );
  NR2SVTX2 U902 ( .A(n163), .B(n164), .Z(n1385) );
  NR2ASVTX2 U903 ( .A(n1220), .B(n974), .Z(n1234) );
  AO7SVTX1 U904 ( .A(n1238), .B(n1232), .C(n1231), .Z(n1233) );
  AO8SVTX1 U905 ( .A(n1356), .B(n1355), .C(n1637), .D(n1354), .Z(n1357) );
  F_IVSVTX0H U906 ( .A(n986), .Z(n1340) );
  AO6SVTX1 U907 ( .A(n988), .B(n985), .C(n1340), .Z(n987) );
  CTIVSVTX4 U908 ( .A(n1253), .Z(n1150) );
  F_AO2SVTX1 U909 ( .A(n1296), .B(n1533), .C(n65), .D(n1532), .Z(n1534) );
  F_AO2SVTX1 U910 ( .A(n1596), .B(n1554), .C(n65), .D(n1553), .Z(n1555) );
  ENSVTX0H U911 ( .A(n1609), .B(n1608), .Z(n1630) );
  AO1SVTX2 U912 ( .A(n1296), .B(n1204), .C(n1203), .D(n1202), .Z(n1205) );
  AO7ABSVTX4 U913 ( .A(n1596), .B(n325), .C(n324), .Z(m2[14]) );
  AO6SVTX2 U914 ( .A(n4), .B(n323), .C(n322), .Z(n324) );
  NR2SVTX2 U915 ( .A(n1258), .B(n1257), .Z(n44) );
  CTIVSVTX2 U916 ( .A(n579), .Z(n580) );
  AN2SVTX4 U917 ( .A(n1548), .B(n936), .Z(n74) );
  F_AN2SVTX2 U918 ( .A(n632), .B(n630), .Z(n24) );
  F_AN2SVTX2 U919 ( .A(n628), .B(n1065), .Z(n25) );
  ND2SVTX2 U920 ( .A(n125), .B(n230), .Z(n94) );
  NR3ASVTX4 U921 ( .A(n1), .B(n663), .C(n1045), .Z(n664) );
  NR2ASVTX4 U922 ( .A(n1045), .B(n1161), .Z(n1163) );
  ND2SVTX2 U923 ( .A(m1[4]), .B(m1[2]), .Z(n1589) );
  IVSVTX12 U924 ( .A(n1454), .Z(n283) );
  ND2SVTX4 U925 ( .A(n781), .B(n780), .Z(n26) );
  F_AN2SVTX2 U926 ( .A(n1049), .B(n674), .Z(n61) );
  F_ND2ASVTX2 U927 ( .A(n272), .B(m1[2]), .Z(n235) );
  ND2SVTX2 U928 ( .A(n500), .B(n1094), .Z(n460) );
  IVSVTX2 U929 ( .A(n249), .Z(n234) );
  AO20CSVTX8 U930 ( .A(n397), .B(n737), .C(n28), .D(n396), .Z(n27) );
  AO1SVTX8 U931 ( .A(n993), .B(n994), .C(n992), .D(n991), .Z(m2[22]) );
  ND2SVTX2 U932 ( .A(n500), .B(n499), .Z(n501) );
  NR3SVTX2 U933 ( .A(m1[23]), .B(n202), .C(n201), .Z(n204) );
  ND3SVTX4 U934 ( .A(n477), .B(n476), .C(n475), .Z(n487) );
  F_IVSVTX0H U935 ( .A(n245), .Z(n246) );
  NR2SVTX4 U936 ( .A(m1[15]), .B(n188), .Z(n29) );
  NR2SVTX4 U937 ( .A(n30), .B(n189), .Z(n190) );
  IVSVTX4 U938 ( .A(n29), .Z(n30) );
  AN4SVTX6 U939 ( .A(n852), .B(n781), .C(n905), .D(n780), .Z(n77) );
  ND2SVTX2 U940 ( .A(n102), .B(n187), .Z(n86) );
  IVSVTX2 U941 ( .A(n627), .Z(n32) );
  NR2SVTX2 U942 ( .A(n651), .B(m1[22]), .Z(n627) );
  NR2ASVTX4 U943 ( .A(n303), .B(n531), .Z(n197) );
  ND3SVTX4 U944 ( .A(n1239), .B(m1[27]), .C(n195), .Z(n196) );
  NR2SVTX4 U945 ( .A(n604), .B(n575), .Z(n576) );
  AN2SVTX8 U946 ( .A(n93), .B(n34), .Z(n65) );
  NR2ASVTX6 U947 ( .A(n666), .B(n693), .Z(n34) );
  ND2SVTX2 U948 ( .A(n293), .B(m1[13]), .Z(n35) );
  IVSVTX4 U949 ( .A(n199), .Z(n123) );
  ND4ABSVTX4 U950 ( .A(n202), .B(n199), .C(n98), .D(n198), .Z(n99) );
  F_ND2ASVTX2 U951 ( .A(m1[14]), .B(n117), .Z(n469) );
  ND2SVTX2 U952 ( .A(m1[25]), .B(m1[26]), .Z(n36) );
  IVSVTX2 U953 ( .A(n36), .Z(n70) );
  AN2SVTX4 U954 ( .A(n948), .B(n1076), .Z(n37) );
  IVSVTX6 U955 ( .A(m1[21]), .Z(n408) );
  IVSVTX4 U956 ( .A(n7), .Z(n38) );
  AO17SVTX1 U957 ( .A(n857), .B(n1119), .C(n858), .D(n859), .Z(n863) );
  NR2ASVTX2 U958 ( .A(n540), .B(n528), .Z(n769) );
  IVSVTX12 U959 ( .A(n413), .Z(n675) );
  ND3ABSVTX6 U960 ( .A(m1[19]), .B(n651), .C(n90), .Z(n199) );
  ND2SVTX4 U961 ( .A(n943), .B(n1076), .Z(n456) );
  OR2SVTX2 U962 ( .A(n905), .B(n850), .Z(n81) );
  EN3SVTX4 U963 ( .A(n433), .B(n675), .C(n271), .Z(n130) );
  EN3SVTX4 U964 ( .A(n408), .B(n271), .C(n463), .Z(n446) );
  OR2SVTX4 U965 ( .A(m1[13]), .B(n5), .Z(n1263) );
  AO7SVTX1 U966 ( .A(n1329), .B(n1328), .C(n1327), .Z(n1334) );
  NR2SVTX2 U967 ( .A(n385), .B(n1348), .Z(n388) );
  ND2SVTX2 U968 ( .A(n534), .B(n262), .Z(n266) );
  IVSVTX4 U969 ( .A(n340), .Z(n51) );
  NR2SVTX2 U970 ( .A(n220), .B(n1184), .Z(n225) );
  ND3SVTX4 U971 ( .A(n358), .B(n357), .C(n356), .Z(n405) );
  AO7NSVTX4 U972 ( .A(n716), .B(n711), .C(n713), .Z(n439) );
  ND2SVTX2 U973 ( .A(n438), .B(n437), .Z(n713) );
  AO7SVTX8 U974 ( .A(n41), .B(n1169), .C(n48), .Z(n1171) );
  ND2ASVTX8 U975 ( .A(n1341), .B(n1343), .Z(n993) );
  IVSVTX0H U976 ( .A(n1265), .Z(n1642) );
  AO7SVTX1 U977 ( .A(n296), .B(n675), .C(m1[16]), .Z(n128) );
  AO7SVTX6 U978 ( .A(n441), .B(n440), .C(n439), .Z(n442) );
  AO1SVTX4 U979 ( .A(n1296), .B(n903), .C(n902), .D(n901), .Z(n918) );
  IVSVTX2 U980 ( .A(n738), .Z(n892) );
  AO7SVTX2 U981 ( .A(n1279), .B(n754), .C(n753), .Z(n759) );
  NR2SVTX2 U982 ( .A(n747), .B(n746), .Z(n755) );
  F_IVSVTX0H U983 ( .A(n1324), .Z(n921) );
  IVSVTX4 U984 ( .A(n1080), .Z(n944) );
  AO21SVTX6 U985 ( .A(n1096), .B(n1081), .C(n1080), .D(n1079), .Z(n1082) );
  AO6CSVTX8 U986 ( .A(n827), .B(n819), .C(n820), .Z(n1080) );
  AO3ABSVTX4 U987 ( .A(n940), .B(n1094), .C(n939), .D(n1), .Z(n942) );
  NR2ASVTX4 U988 ( .A(n611), .B(n949), .Z(n612) );
  NR4SVTX4 U989 ( .A(n1664), .B(n1096), .C(n1095), .D(n949), .Z(n1097) );
  CTIVSVTX2 U990 ( .A(n559), .Z(n560) );
  ND2SVTX4 U991 ( .A(n731), .B(n349), .Z(n850) );
  AO1ABSVTX6 U992 ( .A(n982), .B(n981), .C(n980), .D(n979), .Z(n983) );
  AO6SVTX1 U993 ( .A(n66), .B(m1[24]), .C(n1116), .Z(n1117) );
  ND2SVTX4 U994 ( .A(n1109), .B(n1067), .Z(n265) );
  IVSVTX4 U995 ( .A(n265), .Z(n304) );
  ND2SVTX2 U996 ( .A(n690), .B(n253), .Z(n907) );
  IVSVTX4 U997 ( .A(n587), .Z(n1065) );
  AO4SVTX1 U998 ( .A(n783), .B(n782), .C(n852), .D(n910), .Z(n784) );
  NR3SVTX2 U999 ( .A(n555), .B(n634), .C(n852), .Z(n556) );
  AO6ABSVTX6 U1000 ( .A(n596), .B(n595), .C(n1650), .Z(n69) );
  AO7SVTX1 U1001 ( .A(n771), .B(n770), .C(n527), .Z(n772) );
  NR3SVTX4 U1002 ( .A(n256), .B(n268), .C(n267), .Z(n269) );
  ND3SVTX4 U1003 ( .A(n1125), .B(m1[23]), .C(n955), .Z(n1060) );
  ND3SVTX2 U1004 ( .A(n944), .B(n1075), .C(n1076), .Z(n945) );
  IVSVTX2 U1005 ( .A(n435), .Z(n436) );
  NR2SVTX2 U1006 ( .A(m1[15]), .B(m1[13]), .Z(n1269) );
  F_ND2ASVTX2 U1007 ( .A(m1[13]), .B(m1[16]), .Z(n1277) );
  NR2SVTX0H U1008 ( .A(n1351), .B(n2), .Z(n1358) );
  ND2SVTX2 U1009 ( .A(n799), .B(n822), .Z(n800) );
  IVSVTX4 U1010 ( .A(n1351), .Z(n182) );
  ND2SVTX2 U1011 ( .A(n49), .B(n263), .Z(n260) );
  NR4ABCSVTX6 U1012 ( .A(n408), .B(n683), .C(n271), .D(n422), .Z(n254) );
  OR2SVTX4 U1013 ( .A(n581), .B(n10), .Z(n80) );
  AO7ABSVTX2 U1014 ( .A(n725), .B(n795), .C(n722), .Z(n730) );
  IVSVTX2 U1015 ( .A(n727), .Z(n721) );
  AO7SVTX2 U1016 ( .A(n958), .B(n956), .C(n65), .Z(n982) );
  ND2ASVTX8 U1017 ( .A(n377), .B(n376), .Z(n963) );
  IVSVTX12 U1018 ( .A(m1[18]), .Z(n271) );
  NR3SVTX8 U1019 ( .A(n146), .B(m1[17]), .C(m1[18]), .Z(n92) );
  NR2SVTX2 U1020 ( .A(m1[0]), .B(m1[1]), .Z(n187) );
  IVSVTX2 U1021 ( .A(n1304), .Z(n1305) );
  ND2SVTX2 U1022 ( .A(n471), .B(n478), .Z(n488) );
  F_AO2SVTX1 U1023 ( .A(n566), .B(m1[7]), .C(n65), .D(n1033), .Z(n1034) );
  ND2SVTX2 U1024 ( .A(n651), .B(n566), .Z(n656) );
  ND2SVTX2 U1025 ( .A(n16), .B(n97), .Z(n201) );
  ND2ASVTX8 U1026 ( .A(n296), .B(n416), .Z(n1368) );
  AO17SVTX4 U1027 ( .A(n1166), .B(n1154), .C(n1152), .D(n1153), .Z(n1157) );
  NR2SVTX2 U1028 ( .A(n117), .B(m1[19]), .Z(n747) );
  FAS1SVTX2 U1029 ( .A(m1[2]), .B(n283), .CI(m1[5]), .CO(n152), .Z(n148) );
  AO6SVTX8 U1030 ( .A(n226), .B(n51), .C(n339), .Z(n780) );
  CTIVSVTX2 U1031 ( .A(n1076), .Z(n1081) );
  ND2SVTX4 U1032 ( .A(n107), .B(n1004), .Z(n109) );
  AO7SVTX1 U1033 ( .A(n762), .B(n1093), .C(n5), .Z(n763) );
  NR2SVTX0H U1034 ( .A(m1[27]), .B(n36), .Z(n667) );
  B_ND2SVTX2 U1035 ( .A(n1398), .B(n1214), .Z(n287) );
  ND2SVTX4 U1036 ( .A(n31), .B(n1409), .Z(n1398) );
  ND2SVTX2 U1037 ( .A(n1394), .B(n1208), .Z(n1179) );
  ND2SVTX2 U1038 ( .A(n535), .B(n310), .Z(n311) );
  ND2SVTX4 U1039 ( .A(n58), .B(n64), .Z(n114) );
  ND4SVTX6 U1040 ( .A(n601), .B(n600), .C(n599), .D(n598), .Z(n602) );
  AO7ABSVTX4 U1041 ( .A(n566), .B(n816), .C(n815), .Z(n1329) );
  AO7NSVTX8 U1042 ( .A(n1238), .B(n764), .C(n763), .Z(n765) );
  ND3ABSVTX6 U1043 ( .A(n1329), .B(n1323), .C(n1325), .Z(n834) );
  ND4ABSVTX8 U1044 ( .A(n785), .B(n77), .C(n784), .D(n1491), .Z(n911) );
  ND2SVTX4 U1045 ( .A(n1160), .B(n1040), .Z(n1044) );
  IVSVTX4 U1046 ( .A(n229), .Z(n125) );
  ND3SVTX8 U1047 ( .A(n126), .B(n312), .C(n671), .Z(n127) );
  AO7SVTX1 U1048 ( .A(m1[16]), .B(m1[19]), .C(m1[18]), .Z(n411) );
  ND2SVTX2 U1049 ( .A(n1162), .B(n1161), .Z(n1337) );
  IVSVTX6 U1050 ( .A(n413), .Z(n416) );
  F_ND3SVTX2 U1051 ( .A(n89), .B(n1487), .C(n293), .Z(n189) );
  NR2SVTX2 U1052 ( .A(n662), .B(n1240), .Z(n1241) );
  NR2SVTX2 U1053 ( .A(n915), .B(n914), .Z(n917) );
  AN3SVTX4 U1054 ( .A(n1050), .B(n1134), .C(n963), .Z(n379) );
  NR2ASVTX2 U1055 ( .A(m1[24]), .B(n229), .Z(n100) );
  IVSVTX12 U1056 ( .A(n316), .Z(n433) );
  IVSVTX2 U1057 ( .A(n723), .Z(n725) );
  ND2SVTX2 U1058 ( .A(n215), .B(n283), .Z(n1477) );
  ND3SVTX4 U1059 ( .A(n960), .B(n383), .C(n382), .Z(n404) );
  ND2SVTX2 U1060 ( .A(n316), .B(n413), .Z(n468) );
  OR2SVTX4 U1061 ( .A(n675), .B(n651), .Z(n63) );
  AO6SVTX2 U1062 ( .A(n547), .B(n6), .C(n399), .Z(n1114) );
  NR2SVTX2 U1063 ( .A(n1046), .B(n1243), .Z(n1047) );
  NR3SVTX8 U1064 ( .A(n74), .B(n942), .C(n941), .Z(n1161) );
  ND2SVTX4 U1065 ( .A(n217), .B(n1022), .Z(n219) );
  IVSVTX4 U1066 ( .A(n1168), .Z(n1169) );
  ND2SVTX4 U1067 ( .A(n1048), .B(n1168), .Z(n1159) );
  ND2SVTX4 U1068 ( .A(n1244), .B(n1247), .Z(n1343) );
  ND2SVTX2 U1069 ( .A(n1248), .B(n1244), .Z(n1245) );
  AO3SVTX2 U1070 ( .A(n668), .B(m1[24]), .C(n667), .D(n666), .Z(n1113) );
  F_ND2SVTX0H U1071 ( .A(m1[24]), .B(m1[23]), .Z(n1128) );
  AN3SVTX4 U1072 ( .A(m1[24]), .B(n1109), .C(n70), .Z(n207) );
  ND2SVTX4 U1073 ( .A(n1247), .B(n1047), .Z(n1168) );
  IVSVTX4 U1074 ( .A(n148), .Z(n1539) );
  BFSVTX12 U1075 ( .A(m1[14]), .Z(n296) );
  NR2SVTX2 U1076 ( .A(n1545), .B(m1[5]), .Z(n1561) );
  F_ND2ASVTX2 U1077 ( .A(n283), .B(n1545), .Z(n91) );
  ND3SVTX2 U1078 ( .A(n1572), .B(n1545), .C(n238), .Z(n191) );
  IVSVTX2 U1079 ( .A(m1[14]), .Z(n1371) );
  ND3ABSVTX6 U1080 ( .A(n375), .B(n744), .C(n374), .Z(n376) );
  OR2ABSVTX4 U1081 ( .A(m1[5]), .B(m1[2]), .Z(n1584) );
  NR2SVTX2 U1082 ( .A(m1[5]), .B(n86), .Z(n97) );
  F_ND2SVTX0H U1083 ( .A(n1409), .B(m1[5]), .Z(n1468) );
  ND3SVTX4 U1084 ( .A(n833), .B(n832), .C(n831), .Z(n1325) );
  ND2SVTX2 U1085 ( .A(m1[13]), .B(n117), .Z(n1276) );
  ND2SVTX4 U1086 ( .A(n271), .B(n117), .Z(n690) );
  ND2SVTX4 U1087 ( .A(n781), .B(n780), .Z(n760) );
  ND2SVTX4 U1088 ( .A(n1300), .B(n1148), .Z(n1152) );
  FAS1SVTX4 U1089 ( .A(m1[13]), .B(m1[12]), .CI(n277), .CO(n132), .Z(n169) );
  NR2SVTX2 U1090 ( .A(n529), .B(n566), .Z(n817) );
  ND2SVTX4 U1091 ( .A(n1296), .B(n705), .Z(n706) );
  ND2ASVTX8 U1092 ( .A(n743), .B(n232), .Z(n674) );
  NR3SVTX2 U1093 ( .A(m1[16]), .B(n675), .C(n462), .Z(n257) );
  CTIVSVTX2 U1094 ( .A(n479), .Z(n470) );
  NR2ASVTX6 U1095 ( .A(n606), .B(n616), .Z(n985) );
  ND2SVTX2 U1096 ( .A(n469), .B(n468), .Z(n479) );
  AN2BSVTX8 U1097 ( .A(n1138), .B(m1[25]), .Z(n303) );
  EO3SVTX4 U1098 ( .A(m1[16]), .B(n296), .C(n675), .Z(n181) );
  ND2ASVTX1 U1099 ( .A(m1[16]), .B(m1[18]), .Z(n731) );
  AO7NSVTX1 U1100 ( .A(n1138), .B(n1060), .C(n65), .Z(n59) );
  IVSVTX2 U1101 ( .A(m1[26]), .Z(n1239) );
  F_MUX21SVTX1 U1102 ( .A(n1069), .B(n1138), .S(n1068), .Z(n73) );
  AN2SVTX4 U1103 ( .A(n715), .B(n714), .Z(n76) );
  IVSVTX4 U1104 ( .A(n256), .Z(n264) );
  ND4SVTX2 U1105 ( .A(n710), .B(n715), .C(n714), .D(n1639), .Z(n723) );
  AN2SVTX0H U1106 ( .A(n701), .B(n63), .Z(n82) );
  NR2ASVTX6 U1107 ( .A(n986), .B(n985), .Z(n1248) );
  NR2SVTX4 U1108 ( .A(m1[27]), .B(m1[26]), .Z(n535) );
  ND2SVTX2 U1109 ( .A(n1138), .B(n535), .Z(n308) );
  ND2SVTX4 U1110 ( .A(n316), .B(n408), .Z(n87) );
  NR3ABSVTX8 U1111 ( .A(n1274), .B(n92), .C(n91), .Z(n198) );
  IVSVTX2 U1112 ( .A(n201), .Z(n98) );
  ND2SVTX4 U1113 ( .A(n100), .B(n99), .Z(n666) );
  ND2SVTX2 U1114 ( .A(n433), .B(m1[18]), .Z(n386) );
  NR2ASVTX6 U1115 ( .A(n271), .B(n433), .Z(n385) );
  NR2SVTX4 U1116 ( .A(n296), .B(n675), .Z(n1346) );
  NR2SVTX2 U1117 ( .A(m1[7]), .B(n277), .Z(n999) );
  NR2SVTX2 U1118 ( .A(m1[6]), .B(n7), .Z(n1424) );
  NR2SVTX2 U1119 ( .A(n999), .B(n1424), .Z(n107) );
  NR2SVTX2 U1120 ( .A(m1[5]), .B(n285), .Z(n1492) );
  NR2SVTX2 U1121 ( .A(m1[7]), .B(n283), .Z(n1460) );
  NR2SVTX2 U1122 ( .A(n1492), .B(n1460), .Z(n1004) );
  NR2SVTX2 U1123 ( .A(n1581), .B(n1586), .Z(n105) );
  ND2SVTX2 U1124 ( .A(m1[0]), .B(n47), .Z(n1530) );
  NR2SVTX2 U1125 ( .A(m1[1]), .B(n283), .Z(n1526) );
  ND2SVTX2 U1126 ( .A(m1[1]), .B(n283), .Z(n1528) );
  ND2SVTX2 U1127 ( .A(n146), .B(m1[6]), .Z(n1583) );
  AO7SVTX4 U1128 ( .A(n1584), .B(n1581), .C(n1583), .Z(n104) );
  ND2SVTX2 U1129 ( .A(m1[7]), .B(n283), .Z(n1495) );
  ND2SVTX2 U1130 ( .A(m1[6]), .B(n7), .Z(n1426) );
  ND2SVTX2 U1131 ( .A(m1[7]), .B(n277), .Z(n1001) );
  NR2SVTX2 U1132 ( .A(n285), .B(n31), .Z(n1210) );
  OR2SVTX2 U1133 ( .A(n7), .B(m1[12]), .Z(n1208) );
  NR2SVTX2 U1134 ( .A(n114), .B(n1179), .Z(n116) );
  ND2SVTX2 U1135 ( .A(n285), .B(n31), .Z(n1393) );
  ND2SVTX2 U1136 ( .A(n7), .B(m1[12]), .Z(n1209) );
  AO6SVTX2 U1137 ( .A(n1208), .B(n111), .C(n110), .Z(n1178) );
  NR2SVTX2 U1138 ( .A(m1[12]), .B(n433), .Z(n1265) );
  ND2SVTX2 U1139 ( .A(m1[12]), .B(n433), .Z(n1643) );
  IVSVTX2 U1140 ( .A(n1264), .Z(n118) );
  AO6ASVTX4 U1141 ( .A(n1643), .B(n1263), .C(n118), .Z(n389) );
  ND2SVTX2 U1142 ( .A(n296), .B(n675), .Z(n1348) );
  AO7SVTX1 U1143 ( .A(n1346), .B(n1349), .C(n1348), .Z(n121) );
  ENSVTX0H U1144 ( .A(n122), .B(n121), .Z(n325) );
  NR2SVTX4 U1145 ( .A(n229), .B(n301), .Z(n309) );
  IVSVTX2 U1146 ( .A(n309), .Z(n126) );
  NR2ASVTX6 U1147 ( .A(n303), .B(n540), .Z(n671) );
  NR2SVTX4 U1148 ( .A(n131), .B(n130), .Z(n717) );
  NR2ASVTX1 U1149 ( .A(n716), .B(n717), .Z(n186) );
  NR2ASVTX6 U1150 ( .A(n136), .B(n167), .Z(n1607) );
  ND2SVTX4 U1151 ( .A(n710), .B(n1639), .Z(n1260) );
  FAS1SVTX4 U1152 ( .A(n296), .B(m1[12]), .CI(n433), .CO(n179), .Z(n174) );
  NR2SVTX4 U1153 ( .A(n181), .B(n180), .Z(n1351) );
  NR2SVTX4 U1154 ( .A(n1353), .B(n1351), .Z(n714) );
  FAS1SVTX4 U1155 ( .A(m1[6]), .B(n7), .CI(n285), .CO(n161), .Z(n160) );
  NR2SVTX2 U1156 ( .A(n160), .B(n159), .Z(n1419) );
  IVSVTX2 U1157 ( .A(n1419), .Z(n140) );
  ND2SVTX2 U1158 ( .A(n139), .B(n138), .Z(n1421) );
  ND2SVTX4 U1159 ( .A(n166), .B(n141), .Z(n431) );
  ND2SVTX2 U1160 ( .A(n143), .B(n142), .Z(n1567) );
  FAS1SVTX2 U1161 ( .A(m1[7]), .B(n283), .CI(m1[6]), .CO(n158), .Z(n154) );
  NR2SVTX4 U1162 ( .A(n155), .B(n154), .Z(n1446) );
  IVSVTX2 U1163 ( .A(n1446), .Z(n144) );
  ND2SVTX4 U1164 ( .A(n1567), .B(n144), .Z(n428) );
  ND2SVTX2 U1165 ( .A(n1539), .B(n145), .Z(n149) );
  F_ENSVTX2 U1166 ( .A(n1523), .B(n146), .Z(n1531) );
  AO7SVTX1 U1167 ( .A(m1[0]), .B(m1[2]), .C(n146), .Z(n147) );
  F_AN2SVTX2 U1168 ( .A(n235), .B(n147), .Z(n1521) );
  ND2SVTX2 U1169 ( .A(n283), .B(n1531), .Z(n1518) );
  AO7SVTX4 U1170 ( .A(n1519), .B(n1521), .C(n1518), .Z(n1542) );
  NR2ASVTX6 U1171 ( .A(n1538), .B(n1539), .Z(n1541) );
  ND2SVTX2 U1172 ( .A(n151), .B(n150), .Z(n156) );
  ND2SVTX4 U1173 ( .A(n153), .B(n152), .Z(n1568) );
  ND2SVTX4 U1174 ( .A(n155), .B(n154), .Z(n1447) );
  AO7SVTX4 U1175 ( .A(n1568), .B(n1446), .C(n1447), .Z(n426) );
  ND2SVTX2 U1176 ( .A(n158), .B(n157), .Z(n1502) );
  ND2SVTX2 U1177 ( .A(n160), .B(n159), .Z(n1420) );
  AO7SVTX2 U1178 ( .A(n1502), .B(n1419), .C(n1420), .Z(n996) );
  ND2SVTX2 U1179 ( .A(n162), .B(n161), .Z(n1387) );
  ND2SVTX2 U1180 ( .A(n164), .B(n163), .Z(n1386) );
  AO7SVTX2 U1181 ( .A(n1387), .B(n18), .C(n1386), .Z(n165) );
  AO7SVTX4 U1182 ( .A(n431), .B(n1503), .C(n430), .Z(n1637) );
  ND2SVTX4 U1183 ( .A(n168), .B(n167), .Z(n1605) );
  AO6ASVTX8 U1184 ( .A(n1352), .B(n182), .C(n2), .Z(n718) );
  AO7SVTX1 U1185 ( .A(n183), .B(n441), .C(n718), .Z(n184) );
  AO8SVTX1 U1186 ( .A(n1356), .B(n714), .C(n1637), .D(n184), .Z(n185) );
  ENSVTX0H U1187 ( .A(n186), .B(n185), .Z(n323) );
  IVSVTX4 U1188 ( .A(m1[19]), .Z(n342) );
  NR2SVTX2 U1189 ( .A(n422), .B(n253), .Z(n1105) );
  NR2SVTX4 U1190 ( .A(m1[12]), .B(n296), .Z(n1646) );
  ND2SVTX4 U1191 ( .A(n1646), .B(n190), .Z(n193) );
  NR2SVTX2 U1192 ( .A(n7), .B(m1[7]), .Z(n238) );
  ND2ASVTX8 U1193 ( .A(n193), .B(n192), .Z(n531) );
  NR2SVTX2 U1194 ( .A(m1[22]), .B(n690), .Z(n194) );
  NR2SVTX4 U1195 ( .A(n199), .B(n200), .Z(n302) );
  AO6SVTX4 U1196 ( .A(n302), .B(n204), .C(n203), .Z(n327) );
  ND3ABSVTX8 U1197 ( .A(n207), .B(n208), .C(n206), .Z(n1491) );
  ND2SVTX2 U1198 ( .A(n277), .B(n1409), .Z(n1402) );
  ND2SVTX2 U1199 ( .A(n1402), .B(n1222), .Z(n1185) );
  ND2SVTX2 U1200 ( .A(m1[12]), .B(n89), .Z(n1188) );
  NR2SVTX2 U1201 ( .A(m1[6]), .B(n1409), .Z(n1432) );
  NR2SVTX2 U1202 ( .A(m1[7]), .B(n102), .Z(n1018) );
  NR2SVTX2 U1203 ( .A(n1432), .B(n1018), .Z(n217) );
  ND2SVTX2 U1204 ( .A(n47), .B(n1523), .Z(n1511) );
  NR2SVTX2 U1205 ( .A(n47), .B(n1523), .Z(n1510) );
  ND2SVTX2 U1206 ( .A(m1[5]), .B(n1572), .Z(n210) );
  F_ND2ASVTX1 U1207 ( .A(m1[4]), .B(m1[2]), .Z(n1574) );
  ND2SVTX2 U1208 ( .A(m1[5]), .B(n276), .Z(n1476) );
  ND2SVTX2 U1209 ( .A(m1[6]), .B(n1409), .Z(n1433) );
  NR2SVTX2 U1210 ( .A(n277), .B(n1409), .Z(n1223) );
  NR2SVTX2 U1211 ( .A(n31), .B(n38), .Z(n1221) );
  ND2SVTX2 U1212 ( .A(n277), .B(n221), .Z(n1186) );
  AO7SVTX2 U1213 ( .A(n1186), .B(n223), .C(n222), .Z(n224) );
  NR2SVTX4 U1214 ( .A(n225), .B(n224), .Z(n341) );
  NR2SVTX2 U1215 ( .A(n221), .B(m1[14]), .Z(n1286) );
  NR2SVTX2 U1216 ( .A(n1274), .B(m1[15]), .Z(n1283) );
  AO7SVTX1 U1217 ( .A(n331), .B(n1655), .C(n338), .Z(n1361) );
  AO6SVTX1 U1218 ( .A(n1361), .B(n1360), .C(n1359), .Z(n227) );
  ENSVTX0H U1219 ( .A(n228), .B(n227), .Z(n321) );
  NR2ASVTX6 U1220 ( .A(n125), .B(n231), .Z(n668) );
  NR2ASVTX6 U1221 ( .A(n671), .B(n668), .Z(n693) );
  ND2SVTX2 U1222 ( .A(m1[15]), .B(n416), .Z(n480) );
  F_ND2ASVTX2 U1223 ( .A(n285), .B(n89), .Z(n1405) );
  NR2SVTX2 U1224 ( .A(n7), .B(n31), .Z(n248) );
  NR2SVTX2 U1225 ( .A(m1[12]), .B(n277), .Z(n1613) );
  NR2SVTX2 U1226 ( .A(n1613), .B(n67), .Z(n249) );
  NR2SVTX2 U1227 ( .A(n1192), .B(n234), .Z(n471) );
  IVSVTX0H U1228 ( .A(n471), .Z(n250) );
  NR2SVTX2 U1229 ( .A(m1[2]), .B(n283), .Z(n1591) );
  NR2SVTX2 U1230 ( .A(m1[1]), .B(n47), .Z(n236) );
  NR2SVTX2 U1231 ( .A(n245), .B(n1025), .Z(n472) );
  AO6SVTX1 U1232 ( .A(n1028), .B(n241), .C(n240), .Z(n477) );
  ND2SVTX2 U1233 ( .A(m1[6]), .B(n283), .Z(n1482) );
  CTIVSVTX2 U1234 ( .A(n242), .Z(n244) );
  F_ND2SVTX0H U1235 ( .A(m1[7]), .B(m1[5]), .Z(n243) );
  AO7SVTX2 U1236 ( .A(n1482), .B(n244), .C(n243), .Z(n1026) );
  ND2SVTX2 U1237 ( .A(n1026), .B(n246), .Z(n476) );
  AO1CDSVTX4 U1238 ( .A(n1481), .B(n472), .C(n477), .D(n476), .Z(n1407) );
  ND2SVTX2 U1239 ( .A(n285), .B(n277), .Z(n1406) );
  ND2SVTX2 U1240 ( .A(n7), .B(n31), .Z(n247) );
  ND2SVTX2 U1241 ( .A(m1[12]), .B(n277), .Z(n1615) );
  NR2SVTX2 U1242 ( .A(n1646), .B(n1269), .Z(n467) );
  F_ND2ASVTX2 U1243 ( .A(n221), .B(n296), .Z(n1647) );
  AO7SVTX1 U1244 ( .A(n1363), .B(n1365), .C(n1364), .Z(n251) );
  ENSVTX0H U1245 ( .A(n252), .B(n251), .Z(n319) );
  NR3ABSVTX8 U1246 ( .A(n255), .B(n254), .C(n531), .Z(n256) );
  ND2SVTX4 U1247 ( .A(n1109), .B(n303), .Z(n538) );
  ND4SVTX4 U1248 ( .A(n257), .B(n271), .C(n398), .D(n627), .Z(n259) );
  NR2ASVTX6 U1249 ( .A(n534), .B(n302), .Z(n268) );
  NR3ABSVTX8 U1250 ( .A(n300), .B(n266), .C(n268), .Z(n528) );
  NR4ABCSVTX6 U1251 ( .A(n540), .B(n768), .C(n263), .D(n528), .Z(n270) );
  NR2SVTX8 U1252 ( .A(n270), .B(n269), .Z(n578) );
  CTIVSVTX4 U1253 ( .A(n368), .Z(n367) );
  ND2SVTX2 U1254 ( .A(m1[6]), .B(n1572), .Z(n1559) );
  ND2SVTX2 U1255 ( .A(n1523), .B(n283), .Z(n1515) );
  NR2SVTX2 U1256 ( .A(n1523), .B(n283), .Z(n1514) );
  ND2SVTX2 U1257 ( .A(m1[5]), .B(n1545), .Z(n1560) );
  NR2SVTX4 U1258 ( .A(n275), .B(n274), .Z(n292) );
  ND2SVTX4 U1259 ( .A(n38), .B(m1[12]), .Z(n1214) );
  NR2SVTX2 U1260 ( .A(n1409), .B(m1[5]), .Z(n1467) );
  ND2SVTX2 U1261 ( .A(n1458), .B(n278), .Z(n1014) );
  IVSVTX4 U1262 ( .A(n281), .Z(n291) );
  F_ND2ASVTX2 U1263 ( .A(m1[7]), .B(n283), .Z(n1469) );
  AO7SVTX2 U1264 ( .A(n1469), .B(n1467), .C(n1468), .Z(n1012) );
  NR2SVTX2 U1265 ( .A(n7), .B(n215), .Z(n1429) );
  NR2ASVTX6 U1266 ( .A(n285), .B(n31), .Z(n1397) );
  NR2SVTX2 U1267 ( .A(m1[12]), .B(n38), .Z(n1213) );
  ND2SVTX4 U1268 ( .A(n1277), .B(n1652), .Z(n295) );
  ND2SVTX2 U1269 ( .A(m1[13]), .B(n89), .Z(n1619) );
  NR2SVTX2 U1270 ( .A(n89), .B(m1[13]), .Z(n1618) );
  NR2SVTX2 U1271 ( .A(m1[14]), .B(n293), .Z(n1195) );
  AO6SVTX2 U1272 ( .A(n1618), .B(n1196), .C(n1195), .Z(n1278) );
  NR2SVTX2 U1273 ( .A(n221), .B(m1[15]), .Z(n1651) );
  AO6SVTX4 U1274 ( .A(n1620), .B(n373), .C(n748), .Z(n1369) );
  AO7SVTX1 U1275 ( .A(n297), .B(n1369), .C(n1367), .Z(n298) );
  ND3SVTX4 U1276 ( .A(n301), .B(n302), .C(n300), .Z(n307) );
  ND3SVTX2 U1277 ( .A(n303), .B(n305), .C(n304), .Z(n306) );
  NR2SVTX4 U1278 ( .A(n309), .B(n308), .Z(n313) );
  AO6SVTX2 U1279 ( .A(n65), .B(n319), .C(n318), .Z(n320) );
  AO7SVTX2 U1280 ( .A(n1238), .B(n321), .C(n320), .Z(n322) );
  IVSVTX4 U1281 ( .A(n327), .Z(n328) );
  NR2SVTX4 U1282 ( .A(n668), .B(n328), .Z(n669) );
  ND2SVTX4 U1283 ( .A(n329), .B(n669), .Z(n1049) );
  IVSVTX4 U1284 ( .A(n1049), .Z(n529) );
  ND3ABSVTX8 U1285 ( .A(n330), .B(n340), .C(n1403), .Z(n781) );
  ND2SVTX2 U1286 ( .A(n651), .B(n271), .Z(n849) );
  ND2SVTX2 U1287 ( .A(n347), .B(n849), .Z(n555) );
  NR2SVTX2 U1288 ( .A(n552), .B(n634), .Z(n352) );
  NR2SVTX2 U1289 ( .A(n1138), .B(m1[22]), .Z(n1084) );
  AO7SVTX2 U1290 ( .A(n851), .B(n855), .C(n854), .Z(n638) );
  ND2SVTX2 U1291 ( .A(n462), .B(n1139), .Z(n553) );
  AO7SVTX2 U1292 ( .A(n552), .B(n350), .C(n553), .Z(n351) );
  ND2SVTX4 U1293 ( .A(n354), .B(n3), .Z(n357) );
  AO7SVTX2 U1294 ( .A(n926), .B(n928), .C(n925), .Z(n361) );
  ND2SVTX2 U1295 ( .A(n462), .B(n1138), .Z(n961) );
  F_ND2ASVTX2 U1296 ( .A(n416), .B(n651), .Z(n791) );
  ND2SVTX2 U1297 ( .A(n791), .B(n364), .Z(n866) );
  NR2SVTX2 U1298 ( .A(n866), .B(n365), .Z(n1134) );
  ND2SVTX4 U1299 ( .A(n1368), .B(n368), .Z(n752) );
  ND2SVTX4 U1300 ( .A(n371), .B(n370), .Z(n377) );
  NR2SVTX4 U1301 ( .A(n1346), .B(n385), .Z(n390) );
  CTIVSVTX2 U1302 ( .A(n386), .Z(n387) );
  AO3CDSVTX6 U1303 ( .A(n389), .B(n392), .C(n388), .D(n387), .Z(n737) );
  NR2SVTX4 U1304 ( .A(n392), .B(n391), .Z(n738) );
  NR2ASVTX6 U1305 ( .A(n738), .B(n393), .Z(n397) );
  NR2SVTX2 U1306 ( .A(m1[18]), .B(n567), .Z(n889) );
  ND2SVTX2 U1307 ( .A(n735), .B(n63), .Z(n895) );
  ND2SVTX2 U1308 ( .A(n5), .B(m1[19]), .Z(n736) );
  CTIVSVTX2 U1309 ( .A(n736), .Z(n395) );
  ND2SVTX2 U1310 ( .A(n675), .B(n651), .Z(n701) );
  CTIVSVTX2 U1311 ( .A(n701), .Z(n394) );
  ND2SVTX2 U1312 ( .A(m1[18]), .B(n567), .Z(n891) );
  NR2SVTX2 U1313 ( .A(n816), .B(m1[22]), .Z(n621) );
  NR2SVTX2 U1314 ( .A(n621), .B(n618), .Z(n548) );
  F_ND2SVTX0H U1315 ( .A(m1[20]), .B(m1[18]), .Z(n407) );
  AO7SVTX2 U1316 ( .A(m1[20]), .B(m1[18]), .C(n567), .Z(n406) );
  ND2SVTX2 U1317 ( .A(n407), .B(n406), .Z(n449) );
  EN3SVTX4 U1318 ( .A(m1[19]), .B(n408), .C(n534), .Z(n448) );
  ND2SVTX4 U1319 ( .A(n410), .B(n409), .Z(n819) );
  F_ND2SVTX0H U1320 ( .A(m1[16]), .B(m1[19]), .Z(n412) );
  ND2SVTX2 U1321 ( .A(n412), .B(n411), .Z(n445) );
  IVSVTX2 U1322 ( .A(n445), .Z(n415) );
  ND2SVTX2 U1323 ( .A(n415), .B(n414), .Z(n881) );
  NR2ASVTX6 U1324 ( .A(n417), .B(n446), .Z(n879) );
  ND2SVTX4 U1325 ( .A(n881), .B(n418), .Z(n826) );
  ND2SVTX2 U1326 ( .A(n421), .B(n420), .Z(n943) );
  NR2SVTX2 U1327 ( .A(n568), .B(n454), .Z(n1076) );
  IVSVTX2 U1328 ( .A(n456), .Z(n425) );
  ND2SVTX2 U1329 ( .A(n948), .B(n425), .Z(n461) );
  IVSVTX2 U1330 ( .A(n461), .Z(n459) );
  IVSVTX2 U1331 ( .A(n426), .Z(n427) );
  AO7SVTX8 U1332 ( .A(n432), .B(n431), .C(n430), .Z(n795) );
  ND2SVTX2 U1333 ( .A(n386), .B(n434), .Z(n437) );
  EN3SVTX4 U1334 ( .A(n271), .B(n5), .C(m1[19]), .Z(n438) );
  NR2SVTX4 U1335 ( .A(n437), .B(n438), .Z(n711) );
  NR2SVTX4 U1336 ( .A(n711), .B(n717), .Z(n435) );
  ND2SVTX4 U1337 ( .A(n714), .B(n435), .Z(n440) );
  NR2SVTX4 U1338 ( .A(n1260), .B(n440), .Z(n796) );
  NR2SVTX4 U1339 ( .A(n718), .B(n436), .Z(n443) );
  IVSVTX4 U1340 ( .A(n720), .Z(n441) );
  NR2SVTX8 U1341 ( .A(n443), .B(n442), .Z(n822) );
  ND2SVTX8 U1342 ( .A(n657), .B(n822), .Z(n1094) );
  ND2SVTX2 U1343 ( .A(n449), .B(n448), .Z(n820) );
  ND2SVTX2 U1344 ( .A(n943), .B(n1078), .Z(n455) );
  IVSVTX2 U1345 ( .A(n499), .Z(n457) );
  NR2SVTX2 U1346 ( .A(n567), .B(n1136), .Z(n584) );
  NR2SVTX2 U1347 ( .A(n584), .B(n627), .Z(n493) );
  IVSVTX2 U1348 ( .A(n493), .Z(n1066) );
  F_IVSVTX1 U1349 ( .A(n907), .Z(n466) );
  NR2SVTX2 U1350 ( .A(m1[19]), .B(n462), .Z(n838) );
  CTIVSVTX2 U1351 ( .A(n838), .Z(n464) );
  ND2SVTX2 U1352 ( .A(n464), .B(n835), .Z(n492) );
  NR2SVTX2 U1353 ( .A(n1066), .B(n629), .Z(n1125) );
  ND2SVTX2 U1354 ( .A(n416), .B(m1[19]), .Z(n681) );
  ND2SVTX2 U1355 ( .A(n5), .B(m1[18]), .Z(n694) );
  NR2SVTX2 U1356 ( .A(n694), .B(n683), .Z(n490) );
  AO7NSVTX4 U1357 ( .A(n839), .B(n838), .C(n836), .Z(n491) );
  AO17SVTX2 U1358 ( .A(n1125), .B(n691), .C(n494), .D(n65), .Z(n503) );
  F_ND2ASVTX2 U1359 ( .A(n1067), .B(n567), .Z(n586) );
  AO7SVTX1 U1360 ( .A(n584), .B(n625), .C(n586), .Z(n1063) );
  NR2SVTX2 U1361 ( .A(n505), .B(n504), .Z(n508) );
  IVSVTX4 U1362 ( .A(n506), .Z(n507) );
  NR2SVTX4 U1363 ( .A(n1254), .B(n509), .Z(n1041) );
  F_ENSVTX2 U1364 ( .A(n510), .B(n514), .Z(n515) );
  ND2SVTX4 U1365 ( .A(n1596), .B(n515), .Z(n525) );
  ND2SVTX4 U1366 ( .A(n781), .B(n780), .Z(n1119) );
  ND2SVTX2 U1367 ( .A(n26), .B(n1118), .Z(n518) );
  IVSVTX2 U1368 ( .A(n1118), .Z(n520) );
  ND2SVTX4 U1369 ( .A(n522), .B(n521), .Z(n523) );
  ND2SVTX4 U1370 ( .A(n954), .B(n525), .Z(n526) );
  F_ND2SVTX0H U1371 ( .A(m1[25]), .B(m1[24]), .Z(n536) );
  AO7SVTX2 U1372 ( .A(n1106), .B(n541), .C(n540), .Z(n542) );
  ENSVTX4 U1373 ( .A(n550), .B(n549), .Z(n551) );
  CTIVSVTX2 U1374 ( .A(n634), .Z(n561) );
  ND4SVTX2 U1375 ( .A(n345), .B(n562), .C(n561), .D(n1119), .Z(n563) );
  ND4SVTX4 U1376 ( .A(n563), .B(n1491), .C(n564), .D(n565), .Z(n601) );
  CTIVSVTX2 U1377 ( .A(n820), .Z(n572) );
  NR2SVTX2 U1378 ( .A(n569), .B(n568), .Z(n570) );
  ND2SVTX4 U1379 ( .A(n827), .B(n570), .Z(n571) );
  NR2ASVTX6 U1380 ( .A(n653), .B(n609), .Z(n575) );
  NR2SVTX4 U1381 ( .A(n576), .B(n577), .Z(n600) );
  ND2ASVTX6 U1382 ( .A(n1135), .B(n963), .Z(n579) );
  ND2ASVTX4 U1383 ( .A(n581), .B(n580), .Z(n582) );
  ND4SVTX6 U1384 ( .A(n960), .B(n80), .C(n583), .D(n582), .Z(n599) );
  ND2SVTX2 U1385 ( .A(n586), .B(n585), .Z(n596) );
  CTIVSVTX2 U1386 ( .A(n596), .Z(n588) );
  NR2SVTX2 U1387 ( .A(n588), .B(n591), .Z(n589) );
  ND2SVTX4 U1388 ( .A(n589), .B(n595), .Z(n590) );
  IVSVTX4 U1389 ( .A(n590), .Z(n594) );
  NR2SVTX2 U1390 ( .A(n596), .B(n592), .Z(n593) );
  NR2SVTX6 U1391 ( .A(n603), .B(n602), .Z(n616) );
  NR2SVTX2 U1392 ( .A(n989), .B(n1243), .Z(n994) );
  NR2ASVTX2 U1393 ( .A(n652), .B(n937), .Z(n611) );
  ND2SVTX4 U1394 ( .A(n608), .B(n607), .Z(n615) );
  NR2SVTX4 U1395 ( .A(n615), .B(n614), .Z(n617) );
  ND2SVTX4 U1396 ( .A(n617), .B(n616), .Z(n1160) );
  F_ENSVTX2 U1397 ( .A(n84), .B(n623), .Z(n624) );
  NR2SVTX2 U1398 ( .A(n33), .B(n626), .Z(n632) );
  CTIVSVTX2 U1399 ( .A(n629), .Z(n630) );
  NR2SVTX0H U1400 ( .A(n632), .B(n630), .Z(n631) );
  ND2SVTX2 U1401 ( .A(n65), .B(n633), .Z(n647) );
  NR2SVTX2 U1402 ( .A(n635), .B(n634), .Z(n642) );
  B_ND2SVTX1 U1403 ( .A(n345), .B(n643), .Z(n644) );
  ND2SVTX4 U1404 ( .A(n650), .B(n649), .Z(n941) );
  IVSVTX4 U1405 ( .A(n657), .Z(n659) );
  IVSVTX4 U1406 ( .A(n822), .Z(n658) );
  AO7SVTX6 U1407 ( .A(n659), .B(n658), .C(n948), .Z(n660) );
  IVSVTX2 U1408 ( .A(n939), .Z(n663) );
  ND2SVTX4 U1409 ( .A(n664), .B(n665), .Z(n1040) );
  IVSVTX2 U1410 ( .A(n669), .Z(n670) );
  NR2ASVTX2 U1411 ( .A(n675), .B(n779), .Z(n680) );
  F_ENSVTX2 U1412 ( .A(n62), .B(n963), .Z(n678) );
  NR2SVTX2 U1413 ( .A(n683), .B(n682), .Z(n695) );
  NR2ASVTX1 U1414 ( .A(n731), .B(n695), .Z(n684) );
  F_MUX21NSVTX1 U1415 ( .A(n685), .B(n731), .S(n695), .Z(n687) );
  NR3ABSVTX2 U1416 ( .A(n685), .B(n695), .C(n26), .Z(n686) );
  ND3SVTX6 U1417 ( .A(n708), .B(n707), .C(n706), .Z(n777) );
  ND2SVTX4 U1418 ( .A(n1319), .B(n709), .Z(n776) );
  ND2SVTX2 U1419 ( .A(n713), .B(n712), .Z(n726) );
  AO6SVTX6 U1420 ( .A(n720), .B(n76), .C(n719), .Z(n727) );
  NR2ASVTX2 U1421 ( .A(n726), .B(n721), .Z(n722) );
  AO7SVTX2 U1422 ( .A(n727), .B(n726), .C(n4), .Z(n728) );
  AN3CSVTX6 U1423 ( .A(n730), .B(n729), .C(n728), .Z(n1303) );
  NR2SVTX2 U1424 ( .A(n733), .B(n732), .Z(n761) );
  AO6SVTX2 U1425 ( .A(n1644), .B(n738), .C(n737), .Z(n739) );
  ND3ABSVTX2 U1426 ( .A(n743), .B(n742), .C(n741), .Z(n767) );
  NR2SVTX2 U1427 ( .A(n752), .B(n744), .Z(n757) );
  NR2SVTX2 U1428 ( .A(n755), .B(n756), .Z(n753) );
  ND3SVTX4 U1429 ( .A(n759), .B(n758), .C(n1548), .Z(n766) );
  ND3ABSVTX4 U1430 ( .A(n773), .B(n772), .C(n817), .Z(n1317) );
  IVSVTX4 U1431 ( .A(n774), .Z(n775) );
  ND2SVTX4 U1432 ( .A(n776), .B(n775), .Z(n809) );
  NR2ASVTX6 U1433 ( .A(m1[18]), .B(n779), .Z(n902) );
  ND2SVTX4 U1434 ( .A(n839), .B(n835), .Z(n910) );
  IVSVTX4 U1435 ( .A(n911), .Z(n786) );
  NR2SVTX4 U1436 ( .A(n902), .B(n786), .Z(n1309) );
  NR2SVTX4 U1437 ( .A(n1308), .B(n1309), .Z(n806) );
  ND2SVTX4 U1438 ( .A(n796), .B(n795), .Z(n821) );
  AN2SVTX4 U1439 ( .A(n822), .B(n821), .Z(n802) );
  NR2SVTX2 U1440 ( .A(n798), .B(n797), .Z(n799) );
  ND2SVTX4 U1441 ( .A(n803), .B(n1314), .Z(n804) );
  F_AN2SVTX2 U1442 ( .A(n811), .B(n810), .Z(n813) );
  ND2SVTX4 U1443 ( .A(n822), .B(n821), .Z(n824) );
  ND3SVTX2 U1444 ( .A(n823), .B(n825), .C(n824), .Z(n833) );
  IVSVTX4 U1445 ( .A(n824), .Z(n880) );
  ND3ABSVTX2 U1446 ( .A(n827), .B(n825), .C(n880), .Z(n832) );
  NR2SVTX2 U1447 ( .A(n1664), .B(n830), .Z(n831) );
  AO17SVTX2 U1448 ( .A(n846), .B(n955), .C(n845), .D(n844), .Z(n847) );
  ND2SVTX4 U1449 ( .A(n848), .B(n83), .Z(n876) );
  NR2SVTX2 U1450 ( .A(n879), .B(n878), .Z(n900) );
  NR2ASVTX2 U1451 ( .A(n882), .B(n883), .Z(n884) );
  IVSVTX4 U1452 ( .A(n885), .Z(n886) );
  ND2SVTX4 U1453 ( .A(n1313), .B(n1311), .Z(n888) );
  IVSVTX4 U1454 ( .A(n888), .Z(n920) );
  NR2SVTX2 U1455 ( .A(n895), .B(n892), .Z(n897) );
  AO6SVTX2 U1456 ( .A(n897), .B(n1644), .C(n896), .Z(n898) );
  F_EOSVTX2 U1457 ( .A(n899), .B(n898), .Z(n903) );
  AO7ABSVTX2 U1458 ( .A(n905), .B(n904), .C(n65), .Z(n913) );
  IVSVTX4 U1459 ( .A(n919), .Z(n1312) );
  ND2SVTX8 U1460 ( .A(n924), .B(n923), .Z(n1247) );
  AO7SVTX6 U1461 ( .A(n1329), .B(n1324), .C(n1323), .Z(n1327) );
  F_ENSVTX2 U1462 ( .A(n935), .B(n934), .Z(n936) );
  AO7ABSVTX4 U1463 ( .A(n946), .B(n945), .C(n4), .Z(n947) );
  NR2ASVTX6 U1464 ( .A(n37), .B(n949), .Z(n977) );
  ND2SVTX2 U1465 ( .A(n955), .B(n1125), .Z(n956) );
  AO6SVTX2 U1466 ( .A(n968), .B(n970), .C(n971), .Z(n973) );
  NR2ASVTX2 U1467 ( .A(n1076), .B(n1080), .Z(n975) );
  ND2SVTX6 U1468 ( .A(n984), .B(n983), .Z(n988) );
  MUX21NSVTX4 U1469 ( .A(n988), .B(n987), .S(n989), .Z(n992) );
  IVSVTX2 U1470 ( .A(n989), .Z(n990) );
  AO7SVTX1 U1471 ( .A(n995), .B(n1503), .C(n1388), .Z(n997) );
  ENSVTX0H U1472 ( .A(n998), .B(n997), .Z(n1008) );
  IVSVTX0H U1473 ( .A(n999), .Z(n1000) );
  AO7SVTX1 U1474 ( .A(n1424), .B(n1427), .C(n1426), .Z(n1005) );
  ENSVTX0H U1475 ( .A(n1006), .B(n1005), .Z(n1007) );
  AO7NSVTX2 U1476 ( .A(n1011), .B(n1563), .C(n1010), .Z(n1470) );
  AO6SVTX1 U1477 ( .A(n1430), .B(n1015), .C(n1429), .Z(n1016) );
  ENSVTX0H U1478 ( .A(n1017), .B(n1016), .Z(n1037) );
  NR2ASVTX1 U1479 ( .A(n1019), .B(n1018), .Z(n1032) );
  AO6SVTX1 U1480 ( .A(n1023), .B(n1022), .C(n1021), .Z(n1434) );
  AO7SVTX1 U1481 ( .A(n1432), .B(n1434), .C(n1433), .Z(n1024) );
  ENSVTX0H U1482 ( .A(n1032), .B(n1031), .Z(n1033) );
  NR2SVTX4 U1483 ( .A(n1042), .B(n1041), .Z(n1043) );
  IVSVTX2 U1484 ( .A(n1045), .Z(n1162) );
  ND2SVTX2 U1485 ( .A(n1138), .B(n1060), .Z(n1069) );
  AO21SVTX2 U1486 ( .A(n1067), .B(n1066), .C(n1065), .D(n1064), .Z(n1068) );
  AO7SVTX1 U1488 ( .A(n1139), .B(n1114), .C(1'b1), .Z(n1072) );
  AO6SVTX2 U1489 ( .A(n1073), .B(n66), .C(n1072), .Z(n1074) );
  ND2SVTX2 U1490 ( .A(n1078), .B(n1077), .Z(n1079) );
  F_ND2SVTX0H U1491 ( .A(m1[26]), .B(n1138), .Z(n1120) );
  ND2SVTX4 U1492 ( .A(n1149), .B(n1250), .Z(n1166) );
  ND2SVTX4 U1493 ( .A(n1253), .B(n1166), .Z(n1246) );
  IVSVTX0H U1494 ( .A(n1108), .Z(n1110) );
  F_MUX21NSVTX1 U1495 ( .A(n1111), .B(n1110), .S(n1109), .Z(n1112) );
  IVSVTX0H U1496 ( .A(n1128), .Z(n1131) );
  AO17NSVTX2 U1497 ( .A(n1131), .B(n1130), .C(n1129), .D(n65), .Z(n1133) );
  NR2ASVTX1 U1498 ( .A(n1136), .B(n1135), .Z(n1142) );
  AO3SVTX1 U1499 ( .A(n10), .B(n1139), .C(n1138), .D(n1137), .Z(n1141) );
  AO1SVTX2 U1500 ( .A(n1142), .B(n963), .C(m1[25]), .D(n1141), .Z(n1240) );
  ND2SVTX2 U1501 ( .A(n960), .B(n1240), .Z(n1145) );
  AO6SVTX1 U1502 ( .A(m1[25]), .B(n566), .C(n1143), .Z(n1144) );
  ND2SVTX2 U1503 ( .A(n1145), .B(n1144), .Z(n1251) );
  NR2SVTX4 U1504 ( .A(n1246), .B(n1155), .Z(n1158) );
  IVSVTX4 U1505 ( .A(n1151), .Z(n1167) );
  ND2SVTX4 U1506 ( .A(n1150), .B(n1167), .Z(n1154) );
  AO1SVTX8 U1507 ( .A(n1159), .B(n1158), .C(n1157), .D(n1156), .Z(m2[24]) );
  AO6SVTX4 U1508 ( .A(n1339), .B(n1337), .C(n1335), .Z(n1164) );
  ENSVTX4 U1509 ( .A(n1165), .B(n1164), .Z(m2[20]) );
  ENSVTX8 U1510 ( .A(n1172), .B(n1171), .Z(m2[23]) );
  IVSVTX2 U1511 ( .A(n1637), .Z(n1606) );
  AO7SVTX2 U1512 ( .A(n1173), .B(n1606), .C(n1634), .Z(n1174) );
  AO7SVTX1 U1513 ( .A(n1179), .B(n1395), .C(n1178), .Z(n1611) );
  AO6SVTX1 U1514 ( .A(n1611), .B(n58), .C(n1180), .Z(n1181) );
  NR2ASVTX1 U1515 ( .A(n1183), .B(n67), .Z(n1194) );
  IVSVTX0H U1516 ( .A(n1403), .Z(n1224) );
  AO7SVTX1 U1517 ( .A(n1185), .B(n1224), .C(n1184), .Z(n1622) );
  IVSVTX0H U1518 ( .A(n1186), .Z(n1187) );
  AO6SVTX1 U1519 ( .A(n1622), .B(n1188), .C(n1187), .Z(n1189) );
  ENSVTX0H U1520 ( .A(n1194), .B(n1189), .Z(n1190) );
  NR2SVTX2 U1521 ( .A(n1238), .B(n1190), .Z(n1203) );
  NR2ASVTX1 U1522 ( .A(n1196), .B(n1195), .Z(n1198) );
  AO6SVTX1 U1523 ( .A(n1620), .B(n1619), .C(n1618), .Z(n1197) );
  ENSVTX0H U1524 ( .A(n1198), .B(n1197), .Z(n1199) );
  F_AO2SVTX1 U1525 ( .A(n1548), .B(n1199), .C(n31), .D(n566), .Z(n1200) );
  AO7SVTX1 U1526 ( .A(n1201), .B(n45), .C(n1200), .Z(n1202) );
  NR2ASVTX1 U1527 ( .A(n1605), .B(n1607), .Z(n1207) );
  ENSVTX0H U1528 ( .A(n1207), .B(n1637), .Z(n1237) );
  AO7SVTX1 U1529 ( .A(n1210), .B(n1395), .C(n1393), .Z(n1211) );
  ENSVTX0H U1530 ( .A(n1212), .B(n1211), .Z(n1235) );
  NR2ASVTX1 U1531 ( .A(n1214), .B(n1213), .Z(n1219) );
  AO7SVTX1 U1532 ( .A(n1217), .B(n1216), .C(n1215), .Z(n1399) );
  AO6SVTX1 U1533 ( .A(n1399), .B(n1398), .C(n1397), .Z(n1218) );
  ENSVTX0H U1534 ( .A(n1219), .B(n1218), .Z(n1220) );
  NR2ASVTX1 U1535 ( .A(n1222), .B(n1221), .Z(n1229) );
  IVSVTX0H U1536 ( .A(n1402), .Z(n1225) );
  AO7SVTX1 U1537 ( .A(n1225), .B(n1224), .C(n1401), .Z(n1226) );
  ENSVTX0H U1538 ( .A(n1229), .B(n1226), .Z(n1232) );
  IVSVTX0H U1539 ( .A(n1405), .Z(n1227) );
  AO7SVTX1 U1540 ( .A(n1227), .B(n1407), .C(n1406), .Z(n1228) );
  ENSVTX0H U1541 ( .A(n1229), .B(n1228), .Z(n1230) );
  F_AO2SVTX1 U1542 ( .A(n566), .B(n7), .C(n65), .D(n1230), .Z(n1231) );
  AO7SVTX4 U1543 ( .A(n1664), .B(n1237), .C(n1236), .Z(m2[8]) );
  AO6SVTX1 U1544 ( .A(n1644), .B(n1642), .C(n1266), .Z(n1267) );
  EOSVTX0H U1545 ( .A(n1268), .B(n1267), .Z(n1295) );
  NR2ASVTX1 U1546 ( .A(n1270), .B(n1269), .Z(n1273) );
  AO7SVTX1 U1547 ( .A(n1646), .B(n1271), .C(n1647), .Z(n1272) );
  ENSVTX0H U1548 ( .A(n1273), .B(n1272), .Z(n1275) );
  AO4SVTX1 U1549 ( .A(n1275), .B(n45), .C(n39), .D(n1274), .Z(n1294) );
  AO7SVTX1 U1550 ( .A(n1280), .B(n1279), .C(n1278), .Z(n1653) );
  AO6SVTX1 U1551 ( .A(n1653), .B(n1652), .C(n1651), .Z(n1281) );
  ENSVTX0H U1552 ( .A(n1282), .B(n1281), .Z(n1292) );
  NR2ASVTX1 U1553 ( .A(n1284), .B(n1283), .Z(n1290) );
  AO7SVTX1 U1554 ( .A(n1288), .B(n1655), .C(n1287), .Z(n1289) );
  ENSVTX0H U1555 ( .A(n1290), .B(n1289), .Z(n1291) );
  AO4SVTX1 U1556 ( .A(n974), .B(n1292), .C(n1238), .D(n1291), .Z(n1293) );
  AO1SVTX4 U1557 ( .A(n1296), .B(n1295), .C(n1294), .D(n1293), .Z(n1297) );
  AO7SVTX4 U1558 ( .A(n1664), .B(n1298), .C(n1297), .Z(m2[12]) );
  IVSVTX2 U1559 ( .A(n1303), .Z(n1306) );
  NR2ASVTX2 U1560 ( .A(n1330), .B(n1332), .Z(n1322) );
  ND3SVTX2 U1561 ( .A(n1326), .B(n1325), .C(n921), .Z(n1328) );
  ENSVTX4 U1562 ( .A(n1334), .B(n1333), .Z(m2[18]) );
  ND2SVTX2 U1563 ( .A(n1337), .B(n1336), .Z(n1338) );
  NR2ASVTX2 U1564 ( .A(n988), .B(n1340), .Z(n1345) );
  AO7SVTX1 U1565 ( .A(n1353), .B(n441), .C(n1352), .Z(n1354) );
  ENSVTX0H U1566 ( .A(n1358), .B(n1357), .Z(n1378) );
  NR2ASVTX1 U1567 ( .A(n1360), .B(n1359), .Z(n1362) );
  ENSVTX0H U1568 ( .A(n1362), .B(n1361), .Z(n1376) );
  NR2ASVTX1 U1569 ( .A(n1364), .B(n1363), .Z(n1366) );
  ENSVTX0H U1570 ( .A(n1366), .B(n1365), .Z(n1374) );
  ENSVTX0H U1571 ( .A(n1370), .B(n1369), .Z(n1372) );
  AO4SVTX1 U1572 ( .A(n974), .B(n1372), .C(n39), .D(n1371), .Z(n1373) );
  AO6SVTX1 U1573 ( .A(n65), .B(n1374), .C(n1373), .Z(n1375) );
  AO6SVTX2 U1574 ( .A(n4), .B(n1378), .C(n1377), .Z(n1379) );
  AO7ABSVTX2 U1575 ( .A(n1296), .B(n1380), .C(n1379), .Z(m2[13]) );
  F_ND2ASVTX2 U1576 ( .A(n1382), .B(n1381), .Z(n1383) );
  NR2ASVTX1 U1577 ( .A(n1386), .B(n18), .Z(n1392) );
  AO7SVTX1 U1578 ( .A(n1390), .B(n1388), .C(n1387), .Z(n1389) );
  ENSVTX0H U1579 ( .A(n1392), .B(n1391), .Z(n1418) );
  EOSVTX0H U1580 ( .A(n1396), .B(n1395), .Z(n1416) );
  NR2ASVTX1 U1581 ( .A(n1398), .B(n1397), .Z(n1400) );
  ENSVTX0H U1582 ( .A(n1400), .B(n1399), .Z(n1414) );
  ENSVTX0H U1583 ( .A(n1404), .B(n1403), .Z(n1412) );
  ENSVTX0H U1584 ( .A(n1408), .B(n1407), .Z(n1410) );
  AO4SVTX1 U1585 ( .A(n1650), .B(n1410), .C(n39), .D(n1409), .Z(n1411) );
  AO6SVTX1 U1586 ( .A(n1491), .B(n1412), .C(n1411), .Z(n1413) );
  AO7SVTX2 U1587 ( .A(n974), .B(n1414), .C(n1413), .Z(n1415) );
  NR2ASVTX1 U1588 ( .A(n1420), .B(n1419), .Z(n1423) );
  ENSVTX0H U1589 ( .A(n1423), .B(n1422), .Z(n1445) );
  EOSVTX0H U1590 ( .A(n1428), .B(n1427), .Z(n1443) );
  ENSVTX0H U1591 ( .A(n1431), .B(n1430), .Z(n1441) );
  NR2ASVTX1 U1592 ( .A(n1433), .B(n1432), .Z(n1436) );
  ENSVTX0H U1593 ( .A(n1436), .B(n1434), .Z(n1439) );
  ENSVTX0H U1594 ( .A(n1436), .B(n1435), .Z(n1437) );
  AO4SVTX1 U1595 ( .A(n1650), .B(n1437), .C(n39), .D(n215), .Z(n1438) );
  AO6SVTX1 U1596 ( .A(n1491), .B(n1439), .C(n1438), .Z(n1440) );
  AO7SVTX2 U1597 ( .A(n974), .B(n1441), .C(n1440), .Z(n1442) );
  NR2ASVTX1 U1598 ( .A(n1447), .B(n1446), .Z(n1450) );
  IVSVTX0H U1599 ( .A(n1567), .Z(n1448) );
  AO7SVTX1 U1600 ( .A(n1448), .B(n1569), .C(n1568), .Z(n1449) );
  ENSVTX0H U1601 ( .A(n1450), .B(n1449), .Z(n1466) );
  NR2ASVTX1 U1602 ( .A(n1477), .B(n1479), .Z(n1451) );
  ENSVTX0H U1603 ( .A(n1451), .B(n1478), .Z(n1457) );
  NR2ASVTX1 U1604 ( .A(n1482), .B(n1484), .Z(n1453) );
  ENSVTX0H U1605 ( .A(n1453), .B(n1481), .Z(n1455) );
  AO4SVTX1 U1606 ( .A(n45), .B(n1455), .C(n39), .D(n1454), .Z(n1456) );
  AO6SVTX1 U1607 ( .A(n1491), .B(n1457), .C(n1456), .Z(n1465) );
  NR2ASVTX1 U1608 ( .A(n1469), .B(n1471), .Z(n1459) );
  ENSVTX0H U1609 ( .A(n1459), .B(n1470), .Z(n1463) );
  ENSVTX0H U1610 ( .A(n1461), .B(n1498), .Z(n1462) );
  F_AO2SVTX1 U1611 ( .A(n1548), .B(n1463), .C(n1462), .D(n1296), .Z(n1464) );
  NR2ASVTX1 U1612 ( .A(n1468), .B(n1467), .Z(n1473) );
  AO7SVTX1 U1613 ( .A(n1471), .B(n1470), .C(n1469), .Z(n1472) );
  ENSVTX0H U1614 ( .A(n1473), .B(n1472), .Z(n1509) );
  IVSVTX0H U1615 ( .A(n1474), .Z(n1475) );
  AO7SVTX1 U1616 ( .A(n1479), .B(n1478), .C(n1477), .Z(n1480) );
  ENSVTX0H U1617 ( .A(n1486), .B(n1480), .Z(n1490) );
  AO7SVTX1 U1618 ( .A(n1484), .B(n1483), .C(n1482), .Z(n1485) );
  ENSVTX0H U1619 ( .A(n1486), .B(n1485), .Z(n1488) );
  AO4SVTX1 U1620 ( .A(n45), .B(n1488), .C(n39), .D(n1487), .Z(n1489) );
  AO6SVTX1 U1621 ( .A(n1491), .B(n1490), .C(n1489), .Z(n1508) );
  IVSVTX0H U1622 ( .A(n1492), .Z(n1493) );
  AO6SVTX1 U1623 ( .A(n1498), .B(n1497), .C(n1496), .Z(n1499) );
  EOSVTX0H U1624 ( .A(n1500), .B(n1499), .Z(n1506) );
  NR2ASVTX1 U1625 ( .A(n1502), .B(n1501), .Z(n1504) );
  ENSVTX0H U1626 ( .A(n1504), .B(n1503), .Z(n1505) );
  F_AO2SVTX1 U1627 ( .A(n1506), .B(n1596), .C(n4), .D(n1505), .Z(n1507) );
  NR2ASVTX1 U1628 ( .A(n1511), .B(n1510), .Z(n1512) );
  ENSVTX0H U1629 ( .A(n1513), .B(n1512), .Z(n1536) );
  NR2ASVTX1 U1630 ( .A(n1515), .B(n1514), .Z(n1516) );
  ENSVTX0H U1631 ( .A(n1521), .B(n1520), .Z(n1522) );
  AO4SVTX1 U1632 ( .A(n39), .B(n1523), .C(n1522), .D(n1664), .Z(n1524) );
  AO6SVTX1 U1633 ( .A(n1548), .B(n1525), .C(n1524), .Z(n1535) );
  IVSVTX0H U1634 ( .A(n1526), .Z(n1527) );
  EOSVTX0H U1635 ( .A(n1530), .B(n1529), .Z(n1533) );
  ENSVTX0H U1636 ( .A(n1531), .B(n235), .Z(n1532) );
  ENSVTX0H U1637 ( .A(n1552), .B(n1575), .Z(n1557) );
  NR2ASVTX1 U1638 ( .A(n1560), .B(n1561), .Z(n1537) );
  ENSVTX0H U1639 ( .A(n1563), .B(n1537), .Z(n1547) );
  NR2ASVTX1 U1640 ( .A(n1539), .B(n1538), .Z(n1540) );
  NR2SVTX2 U1641 ( .A(n1541), .B(n1540), .Z(n1543) );
  ENSVTX0H U1642 ( .A(n1543), .B(n1542), .Z(n1544) );
  AO4SVTX1 U1643 ( .A(n39), .B(n1545), .C(n1544), .D(n1664), .Z(n1546) );
  AO6SVTX1 U1644 ( .A(n1548), .B(n1547), .C(n1546), .Z(n1556) );
  IVSVTX0H U1645 ( .A(n1586), .Z(n1549) );
  EOSVTX0H U1646 ( .A(n1551), .B(n1585), .Z(n1554) );
  ENSVTX0H U1647 ( .A(n1590), .B(n1552), .Z(n1553) );
  NR2ASVTX1 U1648 ( .A(n1559), .B(n1558), .Z(n1566) );
  IVSVTX0H U1649 ( .A(n1560), .Z(n1564) );
  AO7SVTX1 U1650 ( .A(n1564), .B(n1563), .C(n1562), .Z(n1565) );
  ENSVTX0H U1651 ( .A(n1566), .B(n1565), .Z(n1601) );
  ENSVTX0H U1652 ( .A(n1570), .B(n1569), .Z(n1571) );
  AO4SVTX1 U1653 ( .A(n39), .B(n1572), .C(n1571), .D(n1664), .Z(n1600) );
  IVSVTX0H U1654 ( .A(n1573), .Z(n1576) );
  AO7SVTX1 U1655 ( .A(n1576), .B(n1575), .C(n1574), .Z(n1580) );
  IVSVTX0H U1656 ( .A(n1577), .Z(n1578) );
  ENSVTX0H U1657 ( .A(n1580), .B(n1593), .Z(n1598) );
  AO7SVTX1 U1658 ( .A(n1586), .B(n1585), .C(n1584), .Z(n1587) );
  ENSVTX0H U1659 ( .A(n1588), .B(n1587), .Z(n1595) );
  AO7SVTX1 U1660 ( .A(n1591), .B(n1590), .C(n1589), .Z(n1592) );
  ENSVTX0H U1661 ( .A(n1593), .B(n1592), .Z(n1594) );
  F_AO2SVTX1 U1662 ( .A(n1596), .B(n1595), .C(n65), .D(n1594), .Z(n1597) );
  ENSVTX0H U1663 ( .A(n1612), .B(n1611), .Z(n1628) );
  ENSVTX0H U1664 ( .A(n1623), .B(n1616), .Z(n1617) );
  AO4SVTX1 U1665 ( .A(n45), .B(n1617), .C(n39), .D(n89), .Z(n1627) );
  NR2ASVTX1 U1666 ( .A(n1619), .B(n1618), .Z(n1621) );
  ENSVTX0H U1667 ( .A(n1621), .B(n1620), .Z(n1625) );
  ENSVTX0H U1668 ( .A(n1623), .B(n1622), .Z(n1624) );
  AO4SVTX1 U1669 ( .A(n974), .B(n1625), .C(n1238), .D(n1624), .Z(n1626) );
  IVSVTX0H U1670 ( .A(n1635), .Z(n1638) );
  AO7SVTX1 U1671 ( .A(n1635), .B(n1634), .C(n1633), .Z(n1636) );
  AO8SVTX1 U1672 ( .A(n1639), .B(n1638), .C(n1637), .D(n1636), .Z(n1640) );
  ENSVTX0H U1673 ( .A(n1641), .B(n1640), .Z(n1663) );
  ENSVTX0H U1674 ( .A(n1645), .B(n1644), .Z(n1661) );
  ENSVTX0H U1675 ( .A(n1656), .B(n1648), .Z(n1649) );
  AO4SVTX1 U1676 ( .A(n45), .B(n1649), .C(n39), .D(n221), .Z(n1660) );
  NR2ASVTX1 U1677 ( .A(n1652), .B(n1651), .Z(n1654) );
  ENSVTX0H U1678 ( .A(n1654), .B(n1653), .Z(n1658) );
  ENSVTX0H U1679 ( .A(n1656), .B(n1655), .Z(n1657) );
  AO4SVTX1 U1680 ( .A(n974), .B(n1658), .C(n1238), .D(n1657), .Z(n1659) );
endmodule


module remap_top ( num_i, rslt_o );
  input [31:0] num_i;
  output [31:0] rslt_o;
  wire   n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n618;
  wire   [27:0] keyvalues_m1;

  remap re_map ( .m1({keyvalues_m1[27:12], n216, keyvalues_m1[10:3], n618, 
        keyvalues_m1[1:0]}), .m2(rslt_o[26:0]) );
  IVSVTX0H U200 ( .A(n197), .Z(rslt_o[29]) );
  AO6SVTX6 U201 ( .A(n376), .B(rslt_o[28]), .C(n375), .Z(n491) );
  B_ND2SVTX2 U202 ( .A(n179), .B(n301), .Z(n302) );
  IVSVTX10 U203 ( .A(n173), .Z(keyvalues_m1[5]) );
  AO4SVTX4 U204 ( .A(n176), .B(n518), .C(n589), .D(n611), .Z(n367) );
  AO20DSVTX2 U205 ( .A(n316), .B(n369), .C(n315), .D(n530), .Z(n317) );
  MUX21SVTX4 U206 ( .A(n456), .B(n584), .S(n604), .Z(n173) );
  CTIVSVTX2 U207 ( .A(rslt_o[27]), .Z(n175) );
  AO2ABSVTX4 U208 ( .C(n577), .D(n512), .A(n601), .B(n569), .Z(n467) );
  AO7SVTX4 U209 ( .A(n607), .B(n606), .C(n605), .Z(n608) );
  NR2ASVTX1 U210 ( .A(n537), .B(n362), .Z(n253) );
  ND2ASVTX6 U211 ( .A(n597), .B(n596), .Z(n606) );
  CTIVSVTX2 U212 ( .A(n556), .Z(n559) );
  CTIVSVTX2 U213 ( .A(n176), .Z(n174) );
  NR3SVTX4 U214 ( .A(n495), .B(n377), .C(n604), .Z(keyvalues_m1[0]) );
  B_ND2SVTX2 U215 ( .A(n171), .B(n585), .Z(n586) );
  NR2ASVTX4 U216 ( .A(n577), .B(n488), .Z(n483) );
  AO7SVTX1 U217 ( .A(rslt_o[31]), .B(n421), .C(n252), .Z(n254) );
  NR2ASVTX4 U218 ( .A(n497), .B(n544), .Z(n500) );
  ND2SVTX2 U219 ( .A(n551), .B(n550), .Z(n552) );
  MUX21NSVTX4 U220 ( .A(n454), .B(n486), .S(n196), .Z(n216) );
  AO2SVTX4 U221 ( .A(n532), .B(n531), .C(n530), .D(n529), .Z(n533) );
  MUX21NSVTX6 U222 ( .A(n564), .B(n439), .S(n580), .Z(n457) );
  AO6ASVTX2 U223 ( .A(n172), .B(n502), .C(n297), .Z(n518) );
  AO7ABSVTX4 U224 ( .A(n527), .B(n526), .C(n567), .Z(n534) );
  BFSVTX10 U225 ( .A(n577), .Z(rslt_o[27]) );
  BFSVTX6 U226 ( .A(n567), .Z(n587) );
  IVSVTX4 U227 ( .A(n530), .Z(n176) );
  IVSVTX0H U228 ( .A(n201), .Z(n526) );
  IVSVTX2 U229 ( .A(n585), .Z(n501) );
  IVSVTX0H U230 ( .A(n181), .Z(n182) );
  F_ND2ASVTX2 U231 ( .A(n470), .B(n531), .Z(n459) );
  IVSVTX2 U232 ( .A(n464), .Z(n466) );
  IVSVTX4 U233 ( .A(n567), .Z(n463) );
  IVSVTX0H U234 ( .A(n304), .Z(n181) );
  F_ND2SVTX1 U235 ( .A(n260), .B(n313), .Z(n225) );
  F_ND2ASVTX2 U236 ( .A(n351), .B(n350), .Z(n484) );
  ND3SVTX4 U237 ( .A(n469), .B(n595), .C(n468), .Z(n473) );
  ND2ASVTX4 U238 ( .A(n562), .B(n475), .Z(n550) );
  ND2ASVTX4 U239 ( .A(n425), .B(n424), .Z(n485) );
  IVSVTX4 U240 ( .A(n565), .Z(n195) );
  AO7SVTX2 U241 ( .A(n168), .B(n406), .C(n197), .Z(n603) );
  IVSVTX2 U242 ( .A(n476), .Z(n595) );
  CTIVSVTX4 U243 ( .A(n569), .Z(n171) );
  IVSVTX0H U244 ( .A(n541), .Z(n542) );
  IVSVTX2 U245 ( .A(n592), .Z(n214) );
  B_ND2SVTX2 U246 ( .A(n170), .B(n211), .Z(n548) );
  IVSVTX4 U247 ( .A(n434), .Z(n565) );
  OR2SVTX2 U248 ( .A(n538), .B(n427), .Z(n348) );
  ND3ABSVTX4 U249 ( .A(n539), .B(n495), .C(n494), .Z(n496) );
  BFSVTX4 U250 ( .A(n357), .Z(n358) );
  ND3SVTX2 U251 ( .A(n420), .B(n354), .C(n395), .Z(n349) );
  CTIVSVTX2 U252 ( .A(n427), .Z(n430) );
  IVSVTX8 U253 ( .A(n562), .Z(n494) );
  ND2SVTX2 U254 ( .A(n170), .B(n314), .Z(n590) );
  IVSVTX2 U255 ( .A(n479), .Z(n592) );
  BFSVTX8 U256 ( .A(n537), .Z(n543) );
  IVSVTX0H U257 ( .A(n498), .Z(n538) );
  CTBUFSVTX8 U258 ( .A(n396), .Z(rslt_o[30]) );
  ND3ABSVTX4 U259 ( .A(n400), .B(n395), .C(rslt_o[31]), .Z(n506) );
  AO7SVTX4 U260 ( .A(n421), .B(n410), .C(n364), .Z(n365) );
  AO7ABSVTX2 U261 ( .A(n382), .B(n381), .C(n380), .Z(n211) );
  IVSVTX2 U262 ( .A(rslt_o[31]), .Z(n504) );
  IVSVTX0H U263 ( .A(n191), .Z(n296) );
  CTIVSVTX4 U264 ( .A(n411), .Z(n410) );
  IVSVTX0H U265 ( .A(n345), .Z(n200) );
  IVSVTX0H U266 ( .A(n258), .Z(n186) );
  IVSVTX4 U267 ( .A(n549), .Z(n393) );
  IVSVTX2 U268 ( .A(num_i[3]), .Z(n495) );
  IVSVTX4 U269 ( .A(n396), .Z(n313) );
  IVSVTX0H U270 ( .A(num_i[15]), .Z(n400) );
  OR2SVTX4 U271 ( .A(n303), .B(n435), .Z(n427) );
  AO7ABSVTX2 U272 ( .A(n382), .B(n381), .C(n380), .Z(n479) );
  AO7ABSVTX2 U273 ( .A(n395), .B(num_i[21]), .C(n372), .Z(n374) );
  ND2SVTX4 U274 ( .A(n539), .B(n167), .Z(n359) );
  CTIVSVTX2 U275 ( .A(n332), .Z(n333) );
  ND2ASVTX4 U276 ( .A(n517), .B(n395), .Z(n388) );
  BFSVTX8 U277 ( .A(n401), .Z(rslt_o[31]) );
  IVSVTX4 U278 ( .A(n294), .Z(n502) );
  IVSVTX0H U279 ( .A(n284), .Z(n198) );
  BFSVTX2 U280 ( .A(num_i[4]), .Z(n498) );
  IVSVTX6 U281 ( .A(n378), .Z(n411) );
  NR2ASVTX1 U282 ( .A(num_i[6]), .B(n169), .Z(n386) );
  CTIVSVTX4 U283 ( .A(n341), .Z(n342) );
  ND2SVTX6 U284 ( .A(n267), .B(n327), .Z(n391) );
  IVSVTX0H U285 ( .A(n420), .Z(n379) );
  IVSVTX10 U286 ( .A(n404), .Z(n539) );
  ND3SVTX6 U287 ( .A(n266), .B(n265), .C(n264), .Z(n327) );
  BFSVTX6 U288 ( .A(n217), .Z(n192) );
  F_IVSVTX1 U289 ( .A(n403), .Z(n321) );
  IVSVTX2 U290 ( .A(n268), .Z(n212) );
  CTIVSVTX6 U291 ( .A(n169), .Z(n249) );
  NR2SVTX6 U292 ( .A(n403), .B(n169), .Z(n231) );
  BFSVTX4 U293 ( .A(num_i[28]), .Z(n270) );
  NR3ABSVTX6 U294 ( .A(n237), .B(n236), .C(n235), .Z(n283) );
  F_ND3SVTX2 U295 ( .A(n345), .B(n295), .C(n261), .Z(n262) );
  ND4ASVTX4 U296 ( .A(num_i[10]), .B(n278), .C(n277), .D(n276), .Z(n340) );
  IVSVTX10 U297 ( .A(n230), .Z(n169) );
  IVSVTX2 U298 ( .A(n339), .Z(n187) );
  IVSVTX4 U299 ( .A(num_i[30]), .Z(n268) );
  IVSVTX4 U300 ( .A(n190), .Z(n191) );
  IVSVTX4 U301 ( .A(num_i[25]), .Z(n310) );
  BFSVTX2 U302 ( .A(num_i[9]), .Z(n428) );
  IVSVTX8 U303 ( .A(n319), .Z(n230) );
  IVSVTX2 U304 ( .A(num_i[11]), .Z(n339) );
  IVSVTX2 U305 ( .A(num_i[22]), .Z(n345) );
  IVSVTX4 U306 ( .A(num_i[12]), .Z(n421) );
  IVSVTX2 U307 ( .A(num_i[27]), .Z(n203) );
  IVSVTX4 U308 ( .A(num_i[14]), .Z(n517) );
  IVSVTX4 U309 ( .A(num_i[16]), .Z(n286) );
  IVSVTX2 U310 ( .A(num_i[20]), .Z(n284) );
  IVSVTX2 U311 ( .A(num_i[21]), .Z(n285) );
  NR2SVTX4 U312 ( .A(num_i[31]), .B(num_i[29]), .Z(n239) );
  NR2SVTX6 U313 ( .A(num_i[24]), .B(num_i[25]), .Z(n229) );
  ND2SVTX4 U314 ( .A(n225), .B(n311), .Z(n529) );
  IVSVTX2 U315 ( .A(n189), .Z(n371) );
  ND2SVTX4 U316 ( .A(n359), .B(n414), .Z(n434) );
  IVSVTX0H U317 ( .A(n369), .Z(n493) );
  ND2SVTX2 U318 ( .A(n175), .B(n610), .Z(n614) );
  IVSVTX2 U319 ( .A(n371), .Z(n213) );
  F_MUX21NSVTX1 U320 ( .A(num_i[3]), .B(n498), .S(n434), .Z(n361) );
  MUX21NSVTX4 U321 ( .A(n438), .B(n437), .S(n494), .Z(n456) );
  AN2SVTX0H U322 ( .A(n345), .B(num_i[21]), .Z(n167) );
  AO6ABSVTX4 U323 ( .A(n313), .B(n370), .C(n374), .Z(n458) );
  IVSVTX4 U324 ( .A(num_i[18]), .Z(n172) );
  F_AN2SVTX2 U325 ( .A(n209), .B(n476), .Z(n168) );
  AO7SVTX4 U326 ( .A(rslt_o[27]), .B(n487), .C(n407), .Z(n419) );
  B_ND2SVTX2 U327 ( .A(n358), .B(n515), .Z(n523) );
  OR2SVTX4 U328 ( .A(n464), .B(n416), .Z(n218) );
  ND2SVTX2 U329 ( .A(n507), .B(n506), .Z(n525) );
  IVSVTX10 U330 ( .A(n255), .Z(n537) );
  CTIVSVTX2 U331 ( .A(n442), .Z(n445) );
  ND2SVTX8 U332 ( .A(n614), .B(n613), .Z(keyvalues_m1[22]) );
  AO2ABSVTX4 U333 ( .C(rslt_o[27]), .D(n612), .A(n611), .B(n218), .Z(n613) );
  ND3SVTX6 U334 ( .A(n574), .B(n222), .C(n573), .Z(n610) );
  IVSVTX2 U335 ( .A(n590), .Z(n572) );
  ND2ASVTX6 U336 ( .A(n383), .B(n394), .Z(n487) );
  IVSVTX6 U337 ( .A(n528), .Z(n530) );
  OR2SVTX4 U338 ( .A(n471), .B(n591), .Z(n223) );
  IVSVTX2 U339 ( .A(n525), .Z(n527) );
  MUX21NSVTX6 U340 ( .A(n466), .B(n465), .S(n565), .Z(n601) );
  B_ND2SVTX2 U341 ( .A(n529), .B(n171), .Z(n318) );
  IVSVTX2 U342 ( .A(n594), .Z(n184) );
  NR2ASVTX4 U343 ( .A(n541), .B(n543), .Z(n440) );
  NR2SVTX4 U344 ( .A(n377), .B(n361), .Z(keyvalues_m1[1]) );
  CTIVSVTX2 U345 ( .A(n595), .Z(n183) );
  IVSVTX4 U346 ( .A(n474), .Z(n475) );
  IVSVTX2 U347 ( .A(n415), .Z(n416) );
  IVSVTX4 U348 ( .A(n209), .Z(n470) );
  ND2SVTX2 U349 ( .A(n505), .B(n504), .Z(n507) );
  IVSVTX12 U350 ( .A(n537), .Z(n170) );
  B_ND2SVTX2 U351 ( .A(n498), .B(n397), .Z(n366) );
  IVSVTX6 U352 ( .A(n244), .Z(n396) );
  NR2ASVTX2 U353 ( .A(n420), .B(n427), .Z(n425) );
  ND3ABSVTX8 U354 ( .A(n403), .B(n169), .C(n283), .Z(n341) );
  ND2SVTX6 U355 ( .A(n239), .B(n240), .Z(n194) );
  ND2SVTX6 U356 ( .A(n418), .B(n419), .Z(keyvalues_m1[16]) );
  OR2SVTX4 U357 ( .A(n553), .B(n552), .Z(n554) );
  ND3SVTX6 U358 ( .A(n473), .B(n472), .C(n223), .Z(n488) );
  IVSVTX4 U359 ( .A(n463), .Z(n178) );
  AO6ABSVTX6 U360 ( .A(n183), .B(n184), .C(n593), .Z(n596) );
  MUX21NSVTX4 U361 ( .A(n594), .B(n221), .S(n595), .Z(n394) );
  AO7ABSVTX4 U362 ( .A(n521), .B(n498), .C(n256), .Z(n515) );
  ND2SVTX6 U363 ( .A(n170), .B(n570), .Z(n528) );
  AO7ABSVTX2 U364 ( .A(n430), .B(n201), .C(n305), .Z(n308) );
  ND2SVTX2 U365 ( .A(n429), .B(n445), .Z(n555) );
  ND2SVTX6 U366 ( .A(n414), .B(n333), .Z(n347) );
  B_ND2SVTX2 U367 ( .A(n420), .B(n397), .Z(n362) );
  CTIVSVTX2 U368 ( .A(n447), .Z(n450) );
  ND3SVTX6 U369 ( .A(n389), .B(n388), .C(n387), .Z(n426) );
  B_ND2SVTX2 U370 ( .A(n446), .B(n445), .Z(n452) );
  B_ND2SVTX2 U371 ( .A(num_i[7]), .B(n430), .Z(n431) );
  IVSVTX6 U372 ( .A(n293), .Z(n298) );
  ND3ABSVTX8 U373 ( .A(n492), .B(n385), .C(n231), .Z(n401) );
  NR2ASVTX4 U374 ( .A(n428), .B(n427), .Z(n442) );
  NR2SVTX2 U375 ( .A(num_i[31]), .B(n212), .Z(n377) );
  IVSVTX2 U376 ( .A(n247), .Z(n205) );
  IVSVTX4 U377 ( .A(n323), .Z(n215) );
  BFSVTX2 U378 ( .A(num_i[8]), .Z(n420) );
  NR2SVTX6 U379 ( .A(num_i[23]), .B(num_i[22]), .Z(n228) );
  MUX21NSVTX4 U380 ( .A(n484), .B(n485), .S(n562), .Z(n579) );
  ND2SVTX4 U381 ( .A(num_i[15]), .B(n395), .Z(n224) );
  IVSVTX10 U382 ( .A(n539), .Z(n395) );
  NR3SVTX4 U383 ( .A(n385), .B(n220), .C(n403), .Z(n242) );
  AO21SVTX2 U384 ( .A(n443), .B(n442), .C(n441), .D(n393), .Z(n453) );
  NR2SVTX2 U385 ( .A(n441), .B(n443), .Z(n471) );
  AO4ABSVTX8 U386 ( .C(n483), .D(n482), .A(n585), .B(n174), .Z(
        keyvalues_m1[14]) );
  AO2SVTX4 U387 ( .A(n412), .B(num_i[18]), .C(n411), .D(n191), .Z(n464) );
  ND3SVTX2 U388 ( .A(n397), .B(num_i[6]), .C(n396), .Z(n299) );
  AO6SVTX8 U389 ( .A(n508), .B(n567), .C(n180), .Z(n509) );
  AN3SVTX6 U390 ( .A(n201), .B(n492), .C(rslt_o[28]), .Z(n180) );
  NR2SVTX0H U391 ( .A(n170), .B(n518), .Z(n519) );
  MUX21NSVTX6 U392 ( .A(n598), .B(n606), .S(n604), .Z(n599) );
  AO7SVTX8 U393 ( .A(n577), .B(n576), .C(n575), .Z(keyvalues_m1[21]) );
  AO2ABSVTX4 U394 ( .C(n447), .D(n426), .A(n427), .B(n296), .Z(n474) );
  ND2SVTX4 U395 ( .A(n530), .B(n568), .Z(n462) );
  AO3ABSVTX8 U396 ( .A(n508), .B(n171), .C(n534), .D(n533), .Z(n612) );
  IVSVTX4 U397 ( .A(n458), .Z(n508) );
  IVSVTX8 U398 ( .A(n314), .Z(n357) );
  ND3ASVTX2 U399 ( .A(n495), .B(n397), .C(n396), .Z(n398) );
  NR2ASVTX6 U400 ( .A(n238), .B(n294), .Z(n244) );
  IVSVTX6 U401 ( .A(num_i[9]), .Z(n409) );
  ND2SVTX4 U402 ( .A(num_i[15]), .B(n172), .Z(n259) );
  AO2ASVTX2 U403 ( .C(n186), .D(n395), .A(n339), .B(n411), .Z(n399) );
  OR2SVTX8 U404 ( .A(n569), .B(n589), .Z(n222) );
  MUX21NSVTX6 U405 ( .A(n512), .B(n566), .S(n577), .Z(n513) );
  AO2ABSVTX2 U406 ( .C(n488), .D(n604), .A(n528), .B(n601), .Z(n489) );
  IVSVTX8 U407 ( .A(n194), .Z(n217) );
  ND2SVTX4 U408 ( .A(n177), .B(n178), .Z(n179) );
  IVSVTX2 U409 ( .A(n518), .Z(n177) );
  ND2SVTX2 U410 ( .A(n568), .B(n531), .Z(n301) );
  AO6SVTX6 U411 ( .A(n515), .B(rslt_o[28]), .C(n302), .Z(n490) );
  IVSVTX4 U412 ( .A(n188), .Z(n189) );
  AN4SVTX4 U413 ( .A(num_i[1]), .B(n336), .C(n337), .D(n335), .Z(n207) );
  ND3SVTX2 U414 ( .A(n191), .B(n354), .C(n395), .Z(n350) );
  ND3SVTX4 U415 ( .A(n477), .B(n476), .C(n543), .Z(n551) );
  MUX21NSVTX2 U416 ( .A(n581), .B(n582), .S(n476), .Z(n547) );
  MUX21NSVTX6 U417 ( .A(n578), .B(n219), .S(n196), .Z(keyvalues_m1[8]) );
  AO4SVTX4 U418 ( .A(n410), .B(n409), .C(n539), .D(n408), .Z(n465) );
  AN2BSVTX8 U419 ( .A(n465), .B(n478), .Z(n585) );
  AO3SVTX6 U420 ( .A(n589), .B(n463), .C(n462), .D(n461), .Z(n512) );
  AO4ABSVTX4 U421 ( .C(n501), .D(n611), .A(n171), .B(n588), .Z(n514) );
  ND3ABSVTX4 U422 ( .A(n403), .B(n337), .C(n283), .Z(n238) );
  NR3SVTX6 U423 ( .A(n172), .B(n403), .C(n263), .Z(n257) );
  ND3SVTX4 U424 ( .A(n602), .B(n577), .C(n603), .Z(n407) );
  ND2SVTX4 U425 ( .A(n530), .B(n532), .Z(n602) );
  MUX21NSVTX6 U426 ( .A(n564), .B(n563), .S(n562), .Z(n578) );
  AO7SVTX8 U427 ( .A(n433), .B(n432), .C(n431), .Z(n563) );
  ND4SVTX8 U428 ( .A(n192), .B(n251), .C(n250), .D(n444), .Z(n255) );
  MUX21SVTX8 U429 ( .A(n554), .B(n561), .S(n478), .Z(keyvalues_m1[13]) );
  ND2SVTX4 U430 ( .A(n192), .B(n444), .Z(n447) );
  AO7SVTX4 U431 ( .A(n282), .B(n281), .C(n280), .Z(n291) );
  NR3SVTX2 U432 ( .A(num_i[4]), .B(num_i[5]), .C(n336), .Z(n281) );
  AO7SVTX2 U433 ( .A(n441), .B(n443), .C(n447), .Z(n429) );
  NR2SVTX2 U434 ( .A(n470), .B(n469), .Z(n557) );
  IVSVTX6 U435 ( .A(n170), .Z(n469) );
  AO3CDSVTX6 U436 ( .A(n309), .B(rslt_o[31]), .C(n307), .D(n308), .Z(n376) );
  IVSVTX2 U437 ( .A(n607), .Z(n185) );
  NR3ABSVTX2 U438 ( .A(num_i[3]), .B(n539), .C(n397), .Z(n202) );
  F_ND2ASVTX2 U439 ( .A(n369), .B(n397), .Z(n370) );
  CTIVSVTX4 U440 ( .A(n566), .Z(n576) );
  IVSVTX4 U441 ( .A(n217), .Z(n435) );
  NR2SVTX2 U442 ( .A(num_i[6]), .B(num_i[8]), .Z(n276) );
  IVSVTX2 U443 ( .A(n242), .Z(n243) );
  ND3SVTX1 U444 ( .A(n492), .B(n493), .C(n476), .Z(n497) );
  NR2SVTX2 U445 ( .A(n503), .B(n502), .Z(n505) );
  AO6SVTX1 U446 ( .A(n539), .B(n382), .C(num_i[24]), .Z(n363) );
  NR2SVTX2 U447 ( .A(n405), .B(n404), .Z(n441) );
  BFSVTX0H U448 ( .A(num_i[16]), .Z(n382) );
  IVSVTX2 U449 ( .A(num_i[17]), .Z(n408) );
  AO7SVTX2 U450 ( .A(n422), .B(n397), .C(n384), .Z(n477) );
  B_ND2SVTX0H U451 ( .A(num_i[12]), .B(n169), .Z(n384) );
  NR2SVTX2 U452 ( .A(n170), .B(n390), .Z(n594) );
  IVSVTX2 U453 ( .A(n426), .Z(n390) );
  CTIVSVTX6 U454 ( .A(num_i[10]), .Z(n190) );
  IVSVTX4 U455 ( .A(num_i[7]), .Z(n503) );
  IVSVTX2 U456 ( .A(num_i[24]), .Z(n246) );
  IVSVTX2 U457 ( .A(num_i[19]), .Z(n258) );
  BFSVTX6 U458 ( .A(num_i[17]), .Z(n260) );
  BFSVTX6 U459 ( .A(num_i[23]), .Z(n201) );
  NR2ASVTX1 U460 ( .A(num_i[5]), .B(n539), .Z(n541) );
  IVSVTX4 U461 ( .A(num_i[6]), .Z(n540) );
  F_AN2SVTX2 U462 ( .A(n447), .B(n436), .Z(n437) );
  AN2SVTX0H U463 ( .A(num_i[6]), .B(n404), .Z(n436) );
  AO4SVTX2 U464 ( .A(n427), .B(n495), .C(n503), .D(n356), .Z(n439) );
  NR2ASVTX2 U465 ( .A(n549), .B(n548), .Z(n553) );
  IVSVTX2 U466 ( .A(n555), .Z(n560) );
  NR2SVTX2 U467 ( .A(n592), .B(n591), .Z(n593) );
  CTIVSVTX12 U468 ( .A(n531), .Z(n611) );
  NR2SVTX2 U469 ( .A(num_i[8]), .B(n428), .Z(n280) );
  IVSVTX2 U470 ( .A(num_i[26]), .Z(n295) );
  IVSVTX2 U471 ( .A(num_i[13]), .Z(n188) );
  IVSVTX2 U472 ( .A(n391), .Z(n392) );
  AO2SVTX4 U473 ( .A(n524), .B(n604), .C(n523), .D(n522), .Z(keyvalues_m1[27])
         );
  MUX21NSVTX4 U474 ( .A(n438), .B(n484), .S(n562), .Z(n219) );
  MUX21NSVTX4 U475 ( .A(n555), .B(n563), .S(n494), .Z(n486) );
  MUX21NSVTX4 U476 ( .A(n485), .B(n475), .S(n562), .Z(n454) );
  IVSVTX2 U477 ( .A(n218), .Z(n588) );
  AO7SVTX2 U478 ( .A(num_i[7]), .B(n338), .C(n337), .Z(n344) );
  CTIVSVTX4 U479 ( .A(n170), .Z(n197) );
  OR2SVTX4 U480 ( .A(n379), .B(n378), .Z(n380) );
  ND4SVTX2 U481 ( .A(n249), .B(n403), .C(num_i[6]), .D(n356), .Z(n389) );
  MUX21NSVTX6 U482 ( .A(n440), .B(n439), .S(rslt_o[28]), .Z(n584) );
  AO7ABSVTX8 U483 ( .A(n487), .B(n185), .C(n489), .Z(keyvalues_m1[15]) );
  AO1ASVTX6 U484 ( .A(n453), .B(n452), .C(n451), .D(n556), .Z(n455) );
  MUX21NSVTX4 U485 ( .A(n584), .B(n583), .S(n604), .Z(keyvalues_m1[4]) );
  ND2SVTX4 U486 ( .A(n187), .B(n395), .Z(n449) );
  AO7SVTX4 U487 ( .A(n288), .B(n287), .C(n345), .Z(n289) );
  ND2SVTX4 U488 ( .A(n285), .B(n284), .Z(n288) );
  IVSVTX4 U489 ( .A(n322), .Z(n274) );
  AO3SVTX6 U490 ( .A(n458), .B(n176), .C(n460), .D(n459), .Z(n598) );
  AO21ASVTX8 U491 ( .A(n286), .B(n260), .C(n259), .D(n258), .Z(n266) );
  NR2ASVTX4 U492 ( .A(n213), .B(n539), .Z(n443) );
  AO7ABSVTX4 U493 ( .A(n344), .B(n343), .C(n342), .Z(n346) );
  NR2SVTX4 U494 ( .A(n247), .B(n263), .Z(n303) );
  NR3ABSVTX2 U495 ( .A(n172), .B(n260), .C(n319), .Z(n320) );
  ND3ASVTX2 U496 ( .A(n577), .B(n603), .C(n602), .Z(n605) );
  F_AN2SVTX2 U497 ( .A(n193), .B(n340), .Z(n343) );
  AO7NSVTX4 U498 ( .A(n191), .B(n409), .C(n339), .Z(n193) );
  BFSVTX8 U499 ( .A(n604), .Z(n607) );
  AO6ASVTX2 U500 ( .A(rslt_o[30]), .B(num_i[21]), .C(n312), .Z(n315) );
  IVSVTX12 U501 ( .A(n195), .Z(n196) );
  NR2SVTX2 U502 ( .A(n471), .B(n476), .Z(n406) );
  MUX21NSVTX4 U503 ( .A(n490), .B(n524), .S(n577), .Z(keyvalues_m1[26]) );
  IVSVTX4 U504 ( .A(n202), .Z(n448) );
  MUX21NSVTX6 U505 ( .A(n500), .B(n499), .S(n604), .Z(n618) );
  ND3SVTX2 U506 ( .A(n498), .B(n492), .C(rslt_o[28]), .Z(n499) );
  ND2SVTX4 U507 ( .A(n532), .B(n567), .Z(n460) );
  ND4SVTX2 U508 ( .A(n397), .B(num_i[3]), .C(n313), .D(n182), .Z(n305) );
  ND2SVTX4 U509 ( .A(n171), .B(n568), .Z(n368) );
  MUX21NSVTX2 U510 ( .A(n306), .B(n506), .S(n537), .Z(n307) );
  AO3SVTX4 U511 ( .A(n560), .B(rslt_o[28]), .C(n559), .D(n558), .Z(n561) );
  AO7SVTX6 U512 ( .A(n604), .B(n547), .C(n546), .Z(keyvalues_m1[3]) );
  ND3ABSVTX6 U513 ( .A(n391), .B(n549), .C(n298), .Z(n314) );
  IVSVTX2 U514 ( .A(n295), .Z(n199) );
  ND2SVTX4 U515 ( .A(n232), .B(n233), .Z(n334) );
  AO7SVTX1 U516 ( .A(n385), .B(n403), .C(num_i[5]), .Z(n405) );
  AN3CSVTX6 U517 ( .A(n323), .B(n268), .C(num_i[28]), .Z(n265) );
  ND2SVTX4 U518 ( .A(rslt_o[28]), .B(n557), .Z(n558) );
  IVSVTX8 U519 ( .A(n401), .Z(n397) );
  ND3SVTX8 U520 ( .A(n511), .B(n510), .C(n509), .Z(n566) );
  AO2ABSVTX4 U521 ( .C(n577), .D(n610), .A(n611), .B(n601), .Z(n575) );
  AN2SVTX8 U522 ( .A(n449), .B(n448), .Z(n432) );
  IVSVTX4 U523 ( .A(n203), .Z(n204) );
  ND2SVTX4 U524 ( .A(n207), .B(n342), .Z(n206) );
  NR2SVTX2 U525 ( .A(num_i[29]), .B(num_i[18]), .Z(n234) );
  IVSVTX8 U526 ( .A(n570), .Z(n360) );
  ND3ABSVTX6 U527 ( .A(n391), .B(n549), .C(n298), .Z(n570) );
  ND2SVTX4 U528 ( .A(n224), .B(n402), .Z(n209) );
  ND2SVTX8 U529 ( .A(n503), .B(n540), .Z(n210) );
  ND2SVTX2 U530 ( .A(n503), .B(n540), .Z(n282) );
  NR2SVTX4 U531 ( .A(num_i[30]), .B(num_i[29]), .Z(n226) );
  AN2BSVTX2 U532 ( .A(n397), .B(n396), .Z(n521) );
  ND2SVTX4 U533 ( .A(n214), .B(n531), .Z(n461) );
  AN2SVTX8 U534 ( .A(n537), .B(n357), .Z(n531) );
  AO1CSVTX8 U535 ( .A(n587), .B(n571), .C(n368), .D(n367), .Z(n535) );
  AO4ABSVTX6 U536 ( .C(n433), .D(n355), .A(n430), .B(n493), .Z(n564) );
  AO1CSVTX6 U537 ( .A(n358), .B(n376), .C(n318), .D(n317), .Z(n524) );
  MUX21NSVTX4 U538 ( .A(n579), .B(n578), .S(n196), .Z(keyvalues_m1[9]) );
  MUX21NSVTX6 U539 ( .A(n491), .B(n490), .S(n577), .Z(keyvalues_m1[25]) );
  AO17SVTX4 U540 ( .A(rslt_o[28]), .B(n545), .C(n544), .D(n478), .Z(n546) );
  MUX21NSVTX8 U541 ( .A(n535), .B(n491), .S(rslt_o[27]), .Z(keyvalues_m1[24])
         );
  IVSVTX4 U542 ( .A(num_i[29]), .Z(n323) );
  ND2SVTX4 U543 ( .A(n303), .B(n248), .Z(n250) );
  F_MUX21NSVTX1 U544 ( .A(n187), .B(num_i[7]), .S(n537), .Z(n309) );
  NR2SVTX2 U545 ( .A(n496), .B(n537), .Z(n544) );
  ND2SVTX4 U546 ( .A(n537), .B(n570), .Z(n569) );
  ND2SVTX4 U547 ( .A(n476), .B(n543), .Z(n591) );
  NR2SVTX2 U548 ( .A(n197), .B(n542), .Z(n545) );
  NR2SVTX2 U549 ( .A(n548), .B(rslt_o[28]), .Z(n383) );
  ND3SVTX4 U550 ( .A(n329), .B(n328), .C(n327), .Z(n330) );
  ND3SVTX2 U551 ( .A(n205), .B(num_i[25]), .C(n217), .Z(n328) );
  IVSVTX8 U552 ( .A(n492), .Z(n356) );
  NR3SVTX8 U553 ( .A(num_i[5]), .B(num_i[4]), .C(n210), .Z(n335) );
  IVSVTX12 U554 ( .A(n360), .Z(rslt_o[28]) );
  AO7ABSVTX8 U555 ( .A(n604), .B(n598), .C(n467), .Z(keyvalues_m1[19]) );
  ND3SVTX2 U556 ( .A(n550), .B(n551), .C(n478), .Z(n481) );
  ND3ABSVTX6 U557 ( .A(num_i[16]), .B(num_i[18]), .C(n236), .Z(n385) );
  MUX21NSVTX8 U558 ( .A(n219), .B(n457), .S(n196), .Z(keyvalues_m1[7]) );
  ND2SVTX2 U559 ( .A(n532), .B(n171), .Z(n510) );
  MUX21NSVTX6 U560 ( .A(n486), .B(n579), .S(n196), .Z(keyvalues_m1[10]) );
  NR2SVTX2 U561 ( .A(n385), .B(n220), .Z(n248) );
  NR2SVTX2 U562 ( .A(n385), .B(n334), .Z(n245) );
  IVSVTX2 U563 ( .A(n354), .Z(n433) );
  ND2SVTX2 U564 ( .A(n449), .B(n448), .Z(n468) );
  AN3SVTX6 U565 ( .A(n421), .B(n241), .C(n517), .Z(n220) );
  F_AN2SVTX2 U566 ( .A(n537), .B(n477), .Z(n221) );
  NR2SVTX2 U567 ( .A(n218), .B(n528), .Z(n417) );
  NR2SVTX6 U568 ( .A(num_i[28]), .B(num_i[31]), .Z(n227) );
  ND2SVTX8 U569 ( .A(n227), .B(n226), .Z(n492) );
  NR2SVTX4 U570 ( .A(num_i[19]), .B(num_i[17]), .Z(n236) );
  NR2SVTX6 U571 ( .A(num_i[20]), .B(num_i[21]), .Z(n261) );
  ND2SVTX8 U572 ( .A(n228), .B(n261), .Z(n403) );
  NR2SVTX8 U573 ( .A(num_i[27]), .B(num_i[26]), .Z(n326) );
  ND2SVTX8 U574 ( .A(n326), .B(n229), .Z(n319) );
  NR2SVTX2 U575 ( .A(num_i[9]), .B(num_i[11]), .Z(n233) );
  NR2SVTX2 U576 ( .A(num_i[10]), .B(num_i[8]), .Z(n232) );
  NR2SVTX4 U577 ( .A(n189), .B(num_i[14]), .Z(n237) );
  ND4SVTX4 U578 ( .A(n421), .B(n286), .C(n240), .D(n234), .Z(n235) );
  NR2SVTX6 U579 ( .A(num_i[28]), .B(num_i[30]), .Z(n240) );
  ND2SVTX4 U580 ( .A(n217), .B(n230), .Z(n381) );
  NR2SVTX4 U581 ( .A(num_i[13]), .B(num_i[15]), .Z(n241) );
  ND2ASVTX8 U582 ( .A(n381), .B(n243), .Z(n294) );
  ND2ASVTX8 U583 ( .A(n319), .B(n356), .Z(n404) );
  NR2SVTX4 U584 ( .A(n319), .B(n335), .Z(n304) );
  ND2SVTX4 U585 ( .A(n304), .B(n245), .Z(n251) );
  IVSVTX2 U586 ( .A(n326), .Z(n247) );
  ND2SVTX4 U587 ( .A(n310), .B(n246), .Z(n263) );
  ND2SVTX4 U588 ( .A(n403), .B(n249), .Z(n444) );
  AO6SVTX1 U589 ( .A(n539), .B(n198), .C(n270), .Z(n252) );
  AO1ABSVTX2 U590 ( .A(n363), .B(n255), .C(n254), .D(n253), .Z(n256) );
  ND2ASVTX8 U591 ( .A(n492), .B(n257), .Z(n267) );
  NR2SVTX4 U592 ( .A(n263), .B(n262), .Z(n264) );
  ND2SVTX4 U593 ( .A(n204), .B(n268), .Z(n269) );
  AO21DSVTX8 U594 ( .A(n215), .B(n270), .C(n269), .D(num_i[31]), .Z(n322) );
  ND2SVTX4 U595 ( .A(n199), .B(n217), .Z(n273) );
  NR2SVTX2 U596 ( .A(num_i[24]), .B(num_i[26]), .Z(n271) );
  ND3SVTX4 U597 ( .A(n201), .B(n310), .C(n271), .Z(n272) );
  ND2ASVTX8 U598 ( .A(n272), .B(n217), .Z(n329) );
  ND3SVTX8 U599 ( .A(n274), .B(n273), .C(n329), .Z(n549) );
  NR2SVTX2 U600 ( .A(n191), .B(n187), .Z(n279) );
  NR2SVTX2 U601 ( .A(num_i[4]), .B(num_i[5]), .Z(n278) );
  ND2SVTX4 U602 ( .A(num_i[3]), .B(n409), .Z(n275) );
  IVSVTX4 U603 ( .A(n275), .Z(n277) );
  ND2SVTX4 U604 ( .A(n279), .B(n340), .Z(n292) );
  IVSVTX2 U605 ( .A(num_i[2]), .Z(n336) );
  ND3SVTX4 U606 ( .A(num_i[14]), .B(n286), .C(n408), .Z(n287) );
  ND2SVTX4 U607 ( .A(n289), .B(n230), .Z(n290) );
  AO7NSVTX8 U608 ( .A(n435), .B(n290), .C(n268), .Z(n352) );
  AO17ASVTX8 U609 ( .A(n292), .B(n291), .C(n341), .D(n352), .Z(n293) );
  AO7SVTX2 U610 ( .A(n296), .B(n401), .C(n295), .Z(n297) );
  AN2SVTX8 U611 ( .A(n357), .B(n170), .Z(n567) );
  ND2ASVTX8 U612 ( .A(n404), .B(n401), .Z(n378) );
  AO2SVTX2 U613 ( .A(n411), .B(num_i[14]), .C(n200), .D(n395), .Z(n300) );
  ND2SVTX4 U614 ( .A(n300), .B(n299), .Z(n568) );
  IVSVTX4 U615 ( .A(n314), .Z(n580) );
  AO6SVTX1 U616 ( .A(n186), .B(n502), .C(n204), .Z(n306) );
  AO7NSVTX4 U617 ( .A(n409), .B(rslt_o[31]), .C(n310), .Z(n311) );
  IVSVTX2 U618 ( .A(n521), .Z(n316) );
  IVSVTX2 U619 ( .A(num_i[5]), .Z(n369) );
  AO7SVTX1 U620 ( .A(n371), .B(rslt_o[31]), .C(n323), .Z(n312) );
  ND3SVTX4 U621 ( .A(n321), .B(n356), .C(n320), .Z(n325) );
  AO6ABSVTX2 U622 ( .A(n212), .B(n323), .C(n322), .Z(n324) );
  ND2SVTX4 U623 ( .A(n324), .B(n325), .Z(n331) );
  NR2SVTX8 U624 ( .A(n331), .B(n330), .Z(n414) );
  NR3ABSVTX6 U625 ( .A(n517), .B(n213), .C(n401), .Z(n332) );
  IVSVTX4 U626 ( .A(n334), .Z(n337) );
  NR2SVTX2 U627 ( .A(num_i[6]), .B(n369), .Z(n338) );
  ND3SVTX8 U628 ( .A(n206), .B(n359), .C(n346), .Z(n413) );
  NR2SVTX8 U629 ( .A(n347), .B(n413), .Z(n478) );
  IVSVTX12 U630 ( .A(n478), .Z(n577) );
  ND2SVTX4 U631 ( .A(n192), .B(n444), .Z(n354) );
  ND2SVTX4 U632 ( .A(n349), .B(n348), .Z(n438) );
  NR2SVTX2 U633 ( .A(n540), .B(n427), .Z(n351) );
  IVSVTX4 U634 ( .A(n352), .Z(n353) );
  OR2SVTX8 U635 ( .A(n353), .B(n549), .Z(n562) );
  ND2SVTX2 U636 ( .A(n428), .B(n395), .Z(n355) );
  ND2SVTX2 U637 ( .A(n363), .B(n362), .Z(n571) );
  ND2SVTX2 U638 ( .A(n198), .B(n395), .Z(n364) );
  AO6ASVTX8 U639 ( .A(n366), .B(rslt_o[30]), .C(n365), .Z(n589) );
  F_ND2ASVTX2 U640 ( .A(n371), .B(n411), .Z(n372) );
  AO4ABSVTX6 U641 ( .C(n458), .D(n611), .A(n529), .B(n567), .Z(n375) );
  IVSVTX12 U642 ( .A(n577), .Z(n604) );
  ND2SVTX2 U643 ( .A(n498), .B(n539), .Z(n422) );
  ND3SVTX2 U644 ( .A(n385), .B(n356), .C(n386), .Z(n387) );
  ND2SVTX6 U645 ( .A(n393), .B(n392), .Z(n476) );
  ND2SVTX4 U646 ( .A(n399), .B(n398), .Z(n532) );
  ND3SVTX4 U647 ( .A(num_i[7]), .B(n539), .C(n401), .Z(n402) );
  IVSVTX2 U648 ( .A(n502), .Z(n412) );
  NR2ASVTX6 U649 ( .A(n414), .B(n413), .Z(n415) );
  AO6SVTX2 U650 ( .A(n585), .B(n587), .C(n417), .Z(n418) );
  AO7ABSVTX2 U651 ( .A(n395), .B(num_i[12]), .C(n422), .Z(n423) );
  ND2SVTX4 U652 ( .A(n447), .B(n423), .Z(n424) );
  AN2SVTX0H U653 ( .A(n192), .B(n444), .Z(n446) );
  NR3SVTX6 U654 ( .A(n393), .B(n470), .C(n543), .Z(n451) );
  NR3ABSVTX8 U655 ( .A(n476), .B(n450), .C(n432), .Z(n556) );
  MUX21NSVTX8 U656 ( .A(n455), .B(n454), .S(n196), .Z(keyvalues_m1[12]) );
  MUX21NSVTX8 U657 ( .A(n457), .B(n456), .S(n196), .Z(keyvalues_m1[6]) );
  ND2SVTX4 U658 ( .A(n358), .B(n557), .Z(n472) );
  NR2SVTX2 U659 ( .A(n592), .B(n528), .Z(n480) );
  NR2SVTX4 U660 ( .A(n480), .B(n481), .Z(n482) );
  ND3SVTX2 U661 ( .A(n525), .B(n170), .C(rslt_o[28]), .Z(n511) );
  ND2ASVTX8 U662 ( .A(n514), .B(n513), .Z(keyvalues_m1[20]) );
  AO8SVTX1 U663 ( .A(n192), .B(n200), .C(n249), .D(n212), .Z(n516) );
  AO7SVTX1 U664 ( .A(n517), .B(rslt_o[31]), .C(n516), .Z(n520) );
  AO1SVTX2 U665 ( .A(num_i[6]), .B(n521), .C(n520), .D(n519), .Z(n522) );
  IVSVTX4 U666 ( .A(n612), .Z(n536) );
  MUX21NSVTX8 U667 ( .A(n536), .B(n535), .S(rslt_o[27]), .Z(keyvalues_m1[23])
         );
  NR3SVTX2 U668 ( .A(n539), .B(n538), .C(n537), .Z(n581) );
  NR2ASVTX1 U669 ( .A(n492), .B(n540), .Z(n582) );
  ND2SVTX4 U670 ( .A(n568), .B(n567), .Z(n574) );
  ND2SVTX2 U671 ( .A(n572), .B(n571), .Z(n573) );
  MUX21NSVTX2 U672 ( .A(n582), .B(n581), .S(n360), .Z(n583) );
  AO7ABSVTX4 U673 ( .A(n588), .B(n587), .C(n586), .Z(n600) );
  NR2SVTX4 U674 ( .A(n590), .B(n589), .Z(n597) );
  ND2ASVTX8 U675 ( .A(n600), .B(n599), .Z(keyvalues_m1[18]) );
  NR2SVTX2 U676 ( .A(n463), .B(n601), .Z(n609) );
  ND2ASVTX8 U677 ( .A(n609), .B(n608), .Z(keyvalues_m1[17]) );
endmodule

