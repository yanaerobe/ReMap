
module m_rangemapping ( N, O );
  input [31:0] N;
  output [31:0] O;
  wire   n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918;

  ENSVTX1 U294 ( .A(n800), .B(n799), .Z(O[23]) );
  EOSVTX0H U295 ( .A(n810), .B(n809), .Z(O[20]) );
  ENSVTX0H U296 ( .A(n914), .B(n913), .Z(O[19]) );
  EOSVTX0H U297 ( .A(n815), .B(n814), .Z(O[18]) );
  ENSVTX0H U298 ( .A(n918), .B(n917), .Z(O[21]) );
  IVSVTX0H U299 ( .A(n899), .Z(n792) );
  IVSVTX0H U300 ( .A(n838), .Z(n833) );
  IVSVTX0H U301 ( .A(n811), .Z(n812) );
  IVSVTX0H U302 ( .A(n860), .Z(n878) );
  IVSVTX0H U303 ( .A(n801), .Z(n802) );
  IVSVTX0H U304 ( .A(n806), .Z(n807) );
  IVSVTX0H U305 ( .A(n843), .Z(n874) );
  F_FA1SVTX1 U306 ( .A(n697), .B(n696), .CI(n695), .CO(n694), .Z(n698) );
  IVSVTX0H U307 ( .A(n783), .Z(n696) );
  FA1SVTX2 U308 ( .A(n790), .B(n789), .CI(1'b0), .CO(n791), .Z(n785) );
  F_FA1SVTX1 U309 ( .A(n779), .B(n778), .CI(n777), .CO(n786), .Z(n775) );
  NR2ASVTX1 U310 ( .A(n893), .B(n743), .Z(n778) );
  F_FA1SVTX1 U311 ( .A(n782), .B(n781), .CI(n780), .CO(n695), .Z(n790) );
  AO7SVTX1 U312 ( .A(n892), .B(n784), .C(n783), .Z(n789) );
  F_FA1SVTX1 U313 ( .A(n707), .B(n706), .CI(n705), .CO(n781), .Z(n779) );
  NR2ASVTX1 U314 ( .A(n725), .B(n743), .Z(n766) );
  F_FA1SVTX1 U315 ( .A(n720), .B(n719), .CI(n718), .CO(n769), .Z(n768) );
  HA1SVTX1 U316 ( .A(n700), .B(n699), .CO(n706), .S(n771) );
  NR2ASVTX1 U317 ( .A(n744), .B(n743), .Z(n754) );
  AO7SVTX1 U318 ( .A(n751), .B(n701), .C(n750), .Z(n702) );
  F_FA1SVTX1 U319 ( .A(n710), .B(n709), .CI(n708), .CO(n719), .Z(n760) );
  IVSVTX2 U320 ( .A(n750), .Z(n892) );
  F_FA1SVTX1 U321 ( .A(n749), .B(n748), .CI(n747), .CO(n756), .Z(n734) );
  F_IVSVTX1 U322 ( .A(n714), .Z(n688) );
  AO2NSVTX1 U323 ( .A(n701), .B(n633), .C(n686), .D(n691), .Z(n780) );
  IVSVTX0H U324 ( .A(n631), .Z(n633) );
  AO11NSVTX2 U325 ( .A(n782), .B(n684), .C(n683), .D(n681), .E(n444), .F(n687), 
        .Z(n699) );
  EOSVTX0H U326 ( .A(n697), .B(n638), .Z(n687) );
  EOSVTX0H U327 ( .A(n632), .B(n631), .Z(n686) );
  EOSVTX1 U328 ( .A(n707), .B(n646), .Z(n682) );
  EOSVTX1 U329 ( .A(n782), .B(n635), .Z(n681) );
  IVSVTX0H U330 ( .A(n644), .Z(n645) );
  AO6SVTX1 U331 ( .A(n566), .B(n583), .C(n565), .Z(n567) );
  IVSVTX0H U332 ( .A(n707), .Z(n585) );
  IVSVTX0H U333 ( .A(n782), .Z(n586) );
  EOSVTX1 U334 ( .A(n746), .B(n648), .Z(n666) );
  B_ND2SVTX2 U335 ( .A(n647), .B(n628), .Z(n644) );
  EOSVTX1 U336 ( .A(n749), .B(n551), .Z(n649) );
  AO7SVTX2 U337 ( .A(n583), .B(n618), .C(n584), .Z(n707) );
  AO6SVTX1 U338 ( .A(n583), .B(n582), .C(n581), .Z(n584) );
  AO2ASVTX1 U339 ( .C(n610), .D(n574), .A(n564), .B(O[28]), .Z(n573) );
  IVSVTX0H U340 ( .A(n842), .Z(n521) );
  IVSVTX0H U341 ( .A(n859), .Z(n508) );
  IVSVTX0H U342 ( .A(n855), .Z(n872) );
  IVSVTX0H U343 ( .A(n873), .Z(n516) );
  AO11NSVTX2 U344 ( .A(n432), .B(n704), .C(n691), .D(n437), .E(n444), .F(n443), 
        .Z(n530) );
  IVSVTX2 U345 ( .A(n891), .Z(n684) );
  AO6ABSVTX1 U346 ( .A(n420), .B(n618), .C(n617), .Z(n619) );
  EOSVTX1 U347 ( .A(n531), .B(n440), .Z(n449) );
  IVSVTX0H U348 ( .A(n590), .Z(n423) );
  EOSVTX0H U349 ( .A(n529), .B(n446), .Z(n450) );
  AO6ABSVTX1 U350 ( .A(n420), .B(n623), .C(n622), .Z(n624) );
  IVSVTX0H U351 ( .A(n746), .Z(n609) );
  AO6SVTX1 U352 ( .A(n612), .B(n579), .C(n578), .Z(n618) );
  EOSVTX1 U353 ( .A(n520), .B(n453), .Z(n457) );
  BFSVTX8 U354 ( .A(n444), .Z(n701) );
  AO6NSVTX2 U355 ( .A(n420), .B(n419), .C(n418), .Z(n670) );
  AO11SVTX1 U356 ( .A(n615), .B(n614), .C(n613), .D(n612), .E(n611), .F(n610), 
        .Z(n623) );
  AO7SVTX1 U357 ( .A(O[27]), .B(n321), .C(n280), .Z(n655) );
  OR2SVTX2 U358 ( .A(n632), .B(n752), .Z(n891) );
  CTIVSVTX4 U359 ( .A(n721), .Z(n444) );
  AO11SVTX1 U360 ( .A(n613), .B(n614), .C(n412), .D(n612), .E(n592), .F(n610), 
        .Z(n549) );
  B_ND2SVTX2 U361 ( .A(n752), .B(n692), .Z(n721) );
  AO7CNSVTX4 U362 ( .A(n583), .B(n319), .C(n318), .Z(n752) );
  IVSVTX0H U363 ( .A(n601), .Z(n579) );
  IVSVTX0H U364 ( .A(n616), .Z(n544) );
  AO6ABSVTX1 U365 ( .A(O[28]), .B(n317), .C(n316), .Z(n318) );
  AO6ABSVTX1 U366 ( .A(n543), .B(n542), .C(n541), .Z(n601) );
  IVSVTX0H U367 ( .A(n512), .Z(n361) );
  NR2ASVTX1 U368 ( .A(n326), .B(n324), .Z(n463) );
  NR2ASVTX1 U369 ( .A(N[0]), .B(n417), .Z(n326) );
  F_MUX21NSVTX1 U370 ( .A(N[0]), .B(N[1]), .S(O[27]), .Z(n325) );
  IVSVTX0H U371 ( .A(n398), .Z(n394) );
  IVSVTX0H U372 ( .A(n399), .Z(n371) );
  AO4SVTX1 U373 ( .A(n542), .B(n281), .C(n343), .D(n537), .Z(n597) );
  AO4SVTX1 U374 ( .A(n540), .B(n266), .C(n330), .D(n537), .Z(n267) );
  CTIVSVTX6 U375 ( .A(n420), .Z(O[27]) );
  B_ND2SVTX2 U376 ( .A(n583), .B(n278), .Z(n214) );
  NR2ASVTX2 U377 ( .A(n209), .B(n569), .Z(n598) );
  IVSVTX2 U378 ( .A(n272), .Z(n417) );
  IVSVTX0H U379 ( .A(n363), .Z(n366) );
  AO2ABSVTX1 U380 ( .C(N[7]), .D(n411), .A(n281), .B(n338), .Z(n593) );
  AO2ABSVTX1 U381 ( .C(N[5]), .D(n411), .A(n543), .B(n338), .Z(n370) );
  IVSVTX8 U382 ( .A(n420), .Z(n583) );
  ND2ASVTX4 U383 ( .A(O[29]), .B(O[28]), .Z(n599) );
  IVSVTX2 U384 ( .A(O[29]), .Z(n341) );
  CTIVSVTX6 U385 ( .A(n272), .Z(n420) );
  IVSVTX0H U386 ( .A(N[2]), .Z(n344) );
  IVSVTX0H U387 ( .A(N[3]), .Z(n342) );
  IVSVTX0H U388 ( .A(n346), .Z(n247) );
  AO6SVTX1 U389 ( .A(n244), .B(n243), .C(n242), .Z(n248) );
  AO7SVTX1 U390 ( .A(n308), .B(n261), .C(n249), .Z(n260) );
  IVSVTX0H U391 ( .A(n229), .Z(n250) );
  IVSVTX0H U392 ( .A(N[21]), .Z(n539) );
  IVSVTX2 U393 ( .A(n244), .Z(n263) );
  NR3ABSVTX2 U394 ( .A(n223), .B(n222), .C(n242), .Z(n244) );
  IVSVTX0H U395 ( .A(n700), .Z(n626) );
  IVSVTX0H U396 ( .A(n414), .Z(n546) );
  IVSVTX0H U397 ( .A(N[11]), .Z(n283) );
  AO11SVTX1 U398 ( .A(n611), .B(n614), .C(n592), .D(n612), .E(n613), .F(n610), 
        .Z(n607) );
  AO6ABSVTX1 U399 ( .A(n310), .B(n542), .C(n309), .Z(n591) );
  AO2NSVTX1 U400 ( .A(n326), .B(n354), .C(n598), .D(n332), .Z(n472) );
  AO7SVTX1 U401 ( .A(n607), .B(O[27]), .C(n606), .Z(n710) );
  F_MUX21NSVTX1 U402 ( .A(n356), .B(n349), .S(O[27]), .Z(n352) );
  EOSVTX0H U403 ( .A(n527), .B(n448), .Z(n454) );
  AO11SVTX1 U404 ( .A(n592), .B(n614), .C(n414), .D(n612), .E(n412), .F(n610), 
        .Z(n321) );
  CTIVSVTX6 U405 ( .A(n743), .Z(n777) );
  AO21SVTX1 U406 ( .A(N[6]), .B(n538), .C(n263), .D(n225), .Z(n227) );
  F_ND2SVTX0H U407 ( .A(n477), .B(n476), .Z(n478) );
  AO11NSVTX1 U408 ( .A(n507), .B(n704), .C(n691), .D(n499), .E(n701), .F(n501), 
        .Z(n502) );
  AO7SVTX2 U409 ( .A(O[27]), .B(n401), .C(n390), .Z(n534) );
  IVSVTX0H U410 ( .A(n894), .Z(n693) );
  IVSVTX0H U411 ( .A(n557), .Z(n559) );
  OR2SVTX2 U412 ( .A(n773), .B(n772), .Z(n915) );
  IVSVTX0H U413 ( .A(n883), .Z(n889) );
  F_ND2SVTX0H U414 ( .A(n867), .B(n866), .Z(n871) );
  F_ND2SVTX0H U415 ( .A(n819), .B(n433), .Z(n823) );
  EOSVTX0H U416 ( .A(n906), .B(n905), .Z(O[15]) );
  ENSVTX0H U417 ( .A(n818), .B(n817), .Z(O[17]) );
  IVSVTX0H U418 ( .A(n397), .Z(n211) );
  AO6SVTX6 U419 ( .A(n715), .B(n713), .C(n688), .Z(n724) );
  B_ND2SVTX0H U420 ( .A(n740), .B(n739), .Z(n742) );
  B_ND2SVTX0H U421 ( .A(n727), .B(n726), .Z(n729) );
  NR2SVTX4 U422 ( .A(n700), .B(n699), .Z(n738) );
  CTIVSVTX2 U423 ( .A(n907), .Z(n667) );
  AO7SVTX1 U424 ( .A(n672), .B(n908), .C(n671), .Z(n673) );
  AO11NSVTX4 U425 ( .A(n700), .B(n684), .C(n683), .D(n663), .E(n444), .F(n682), 
        .Z(n708) );
  NR2SVTX4 U426 ( .A(n590), .B(n589), .Z(n647) );
  CTIVSVTX4 U427 ( .A(n891), .Z(n704) );
  F_IVSVTX1 U428 ( .A(n697), .Z(n690) );
  B_ND2SVTX2 U429 ( .A(n405), .B(n404), .Z(n434) );
  AO7SVTX4 U430 ( .A(n417), .B(n573), .C(n572), .Z(n782) );
  AO7SVTX1 U431 ( .A(n417), .B(n549), .C(n416), .Z(n418) );
  F_AO2SVTX1 U432 ( .A(n610), .B(n597), .C(n614), .D(n574), .Z(n575) );
  NR2SVTX1 U433 ( .A(n600), .B(n593), .Z(n269) );
  AO11SVTX2 U434 ( .A(n411), .B(N[12]), .C(n410), .D(N[4]), .E(n209), .F(N[20]), .Z(n580) );
  IVSVTX1 U435 ( .A(n593), .Z(n386) );
  AO4SVTX1 U436 ( .A(n540), .B(n276), .C(n342), .D(n537), .Z(n277) );
  IVSVTX4 U437 ( .A(n209), .Z(n540) );
  B_ND2SVTX2 U438 ( .A(n241), .B(n244), .Z(n251) );
  NR2SVTX1 U439 ( .A(N[14]), .B(n543), .Z(n224) );
  AO7SVTX6 U440 ( .A(n801), .B(n804), .C(n803), .Z(n799) );
  AO6SVTX4 U441 ( .A(n914), .B(n911), .C(n763), .Z(n809) );
  CTIVSVTX4 U442 ( .A(n791), .Z(n794) );
  B_ND2SVTX2 U443 ( .A(n762), .B(n761), .Z(n912) );
  F_IVSVTX1 U444 ( .A(n668), .Z(n674) );
  B_ND2SVTX1 U445 ( .A(n647), .B(n660), .Z(n648) );
  AO7SVTX4 U446 ( .A(n623), .B(n583), .C(n619), .Z(n700) );
  B_ND2SVTX2 U447 ( .A(n328), .B(n327), .Z(n336) );
  CTIVSVTX2 U448 ( .A(n214), .Z(n415) );
  F_ND2ASVTX2 U449 ( .A(n583), .B(n278), .Z(n397) );
  ND2ASVTX6 U450 ( .A(n341), .B(n379), .Z(n600) );
  IVSVTX4 U451 ( .A(n569), .Z(n614) );
  NR2ASVTX4 U452 ( .A(n341), .B(O[28]), .Z(n278) );
  ND2ASVTX4 U453 ( .A(n341), .B(O[28]), .Z(n569) );
  ND2ASVTX4 U454 ( .A(O[29]), .B(n209), .Z(n363) );
  IVSVTX4 U455 ( .A(n338), .Z(n209) );
  IVSVTX4 U456 ( .A(n542), .Z(n411) );
  CTIVSVTX2 U457 ( .A(n251), .Z(n255) );
  CTIVSVTX2 U458 ( .A(N[10]), .Z(n275) );
  AO6SVTX6 U459 ( .A(n917), .B(n915), .C(n774), .Z(n804) );
  AO7SVTX4 U460 ( .A(n806), .B(n809), .C(n808), .Z(n917) );
  B_ND2SVTX2 U461 ( .A(n784), .B(n777), .Z(n783) );
  OR2SVTX8 U462 ( .A(n711), .B(n750), .Z(n743) );
  EOSVTX0H U463 ( .A(n723), .B(n724), .Z(n725) );
  AO6SVTX4 U464 ( .A(n525), .B(n843), .C(n524), .Z(n838) );
  OR2SVTX4 U465 ( .A(n707), .B(n705), .Z(n713) );
  CTIVSVTX2 U466 ( .A(n650), .Z(n651) );
  B_ND2SVTX1 U467 ( .A(n746), .B(n745), .Z(n675) );
  B_ND2SVTX2 U468 ( .A(n660), .B(n645), .Z(n646) );
  OR2SVTX2 U469 ( .A(n697), .B(n636), .Z(n629) );
  CTIVSVTX4 U470 ( .A(n426), .Z(n491) );
  IVSVTX0H U471 ( .A(n658), .Z(n639) );
  CTIVSVTX2 U472 ( .A(n710), .Z(n608) );
  CTIVSVTX2 U473 ( .A(n720), .Z(n640) );
  CTIVSVTX2 U474 ( .A(n670), .Z(n587) );
  AO7SVTX4 U475 ( .A(n396), .B(O[27]), .C(n395), .Z(n529) );
  NR2ASVTX2 U476 ( .A(n603), .B(n602), .Z(n625) );
  CTIVSVTX2 U477 ( .A(n580), .Z(n613) );
  MUX21NSVTX2 U478 ( .A(n365), .B(n358), .S(n379), .Z(n507) );
  MUX21NSVTX2 U479 ( .A(n368), .B(n351), .S(n379), .Z(n512) );
  AO39SVTX2 U480 ( .A(n599), .B(n593), .C(n600), .D(n620), .E(n569), .F(n616), 
        .Z(n419) );
  IVSVTX8 U481 ( .A(O[28]), .Z(n379) );
  CTIVSVTX2 U482 ( .A(n370), .Z(n413) );
  B_ND2SVTX2 U483 ( .A(O[28]), .B(n417), .Z(n376) );
  AO4SVTX2 U484 ( .A(n542), .B(n344), .C(n275), .D(n540), .Z(n393) );
  CTIVSVTX2 U485 ( .A(n320), .Z(n392) );
  AO4SVTX2 U486 ( .A(n542), .B(n342), .C(n283), .D(n540), .Z(n385) );
  AO2ABSVTX2 U487 ( .C(N[1]), .D(n411), .A(n337), .B(n338), .Z(n399) );
  AO2ABSVTX2 U488 ( .C(N[4]), .D(n411), .A(n300), .B(n338), .Z(n320) );
  CTIVSVTX2 U489 ( .A(n257), .Z(n258) );
  AO3CDSVTX6 U490 ( .A(O[31]), .B(n248), .C(n247), .D(n246), .Z(O[29]) );
  AO8SVTX1 U491 ( .A(N[9]), .B(n275), .C(n252), .D(n224), .Z(n225) );
  ND2SVTX6 U492 ( .A(n346), .B(n217), .Z(n261) );
  NR2SVTX1 U493 ( .A(N[30]), .B(n287), .Z(n218) );
  NR4SVTX4 U494 ( .A(N[24]), .B(N[27]), .C(N[26]), .D(N[25]), .Z(n217) );
  CTIVSVTX2 U495 ( .A(N[13]), .Z(n543) );
  CTIVSVTX4 U496 ( .A(N[28]), .Z(n298) );
  B_ND2SVTX2 U497 ( .A(n786), .B(n785), .Z(n798) );
  CTIVSVTX2 U498 ( .A(n698), .Z(n793) );
  IVSVTX2 U499 ( .A(n912), .Z(n763) );
  CTIVSVTX2 U500 ( .A(n916), .Z(n774) );
  OR2SVTX4 U501 ( .A(n762), .B(n761), .Z(n911) );
  B_ND2SVTX2 U502 ( .A(n765), .B(n764), .Z(n808) );
  B_ND2SVTX2 U503 ( .A(n773), .B(n772), .Z(n916) );
  FA1SVTX4 U504 ( .A(n771), .B(n770), .CI(n769), .CO(n776), .Z(n772) );
  IVSVTX4 U505 ( .A(n731), .Z(n711) );
  NR2SVTX6 U506 ( .A(n723), .B(n724), .Z(n689) );
  CTIVSVTX2 U507 ( .A(n727), .Z(n685) );
  CTIVSVTX2 U508 ( .A(n839), .Z(n555) );
  B_ND2SVTX2 U509 ( .A(n853), .B(n872), .Z(n845) );
  B_ND2SVTX2 U510 ( .A(n707), .B(n705), .Z(n714) );
  NR2SVTX4 U511 ( .A(n782), .B(n780), .Z(n723) );
  AO6SVTX2 U512 ( .A(n883), .B(n490), .C(n489), .Z(n860) );
  B_ND2SVTX1 U513 ( .A(n749), .B(n747), .Z(n671) );
  B_ND2SVTX2 U514 ( .A(n670), .B(n669), .Z(n908) );
  AO11NSVTX4 U515 ( .A(n707), .B(n684), .C(n683), .D(n682), .E(n444), .F(n681), 
        .Z(n718) );
  B_ND2SVTX2 U516 ( .A(n459), .B(n458), .Z(n511) );
  B_ND2SVTX2 U517 ( .A(n660), .B(n642), .Z(n643) );
  B_ND2SVTX1 U518 ( .A(n691), .B(n492), .Z(n459) );
  B_ND2SVTX2 U519 ( .A(n423), .B(n660), .Z(n424) );
  NR2SVTX6 U520 ( .A(n426), .B(n408), .Z(n660) );
  ENSVTX0H U521 ( .A(n512), .B(n498), .Z(n501) );
  CTIVSVTX2 U522 ( .A(n647), .Z(n659) );
  F_ND2SVTX1 U523 ( .A(n640), .B(n639), .Z(n641) );
  B_ND2SVTX2 U524 ( .A(n452), .B(n491), .Z(n453) );
  CTIVSVTX2 U525 ( .A(n751), .Z(n784) );
  B_ND2SVTX2 U526 ( .A(n609), .B(n608), .Z(n658) );
  B_ND2SVTX2 U527 ( .A(n422), .B(n421), .Z(n590) );
  F_ND2SVTX1 U528 ( .A(n495), .B(n494), .Z(n496) );
  CTIVSVTX2 U529 ( .A(n749), .Z(n588) );
  B_ND2SVTX2 U530 ( .A(n632), .B(n752), .Z(n893) );
  IVSVTX2 U531 ( .A(n632), .Z(n692) );
  B_ND2SVTX2 U532 ( .A(n383), .B(n382), .Z(n384) );
  B_ND2SVTX2 U533 ( .A(n470), .B(n210), .Z(n335) );
  CTIVSVTX2 U534 ( .A(n529), .Z(n405) );
  CTIVSVTX2 U535 ( .A(n554), .Z(n422) );
  CTIVSVTX2 U536 ( .A(n527), .Z(n383) );
  CTIVSVTX2 U537 ( .A(n520), .Z(n382) );
  CTIVSVTX2 U538 ( .A(n432), .Z(n391) );
  CTIVSVTX2 U539 ( .A(n534), .Z(n428) );
  CTIVSVTX2 U540 ( .A(n486), .Z(n210) );
  AO7SVTX2 U541 ( .A(n323), .B(n583), .C(n322), .Z(n554) );
  B_ND2SVTX2 U542 ( .A(n583), .B(n319), .Z(n312) );
  AO4SVTX2 U543 ( .A(n576), .B(n325), .C(n331), .D(n324), .Z(n477) );
  AO4SVTX2 U544 ( .A(n352), .B(n379), .C(n331), .D(n576), .Z(n488) );
  B_ND2SVTX2 U545 ( .A(n455), .B(n369), .Z(n451) );
  AO7SVTX2 U546 ( .A(n417), .B(n381), .C(n380), .Z(n520) );
  CTIVSVTX2 U547 ( .A(n507), .Z(n495) );
  CTIVSVTX2 U548 ( .A(n514), .Z(n455) );
  CTIVSVTX2 U549 ( .A(n598), .Z(n324) );
  CTIVSVTX2 U550 ( .A(n373), .Z(n374) );
  AO7SVTX2 U551 ( .A(n330), .B(n301), .C(n291), .Z(n574) );
  AO2ABSVTX2 U552 ( .C(N[0]), .D(n411), .A(n339), .B(n338), .Z(n398) );
  ND2ASVTX6 U553 ( .A(O[31]), .B(O[30]), .Z(n537) );
  NR2SVTX2 U554 ( .A(O[31]), .B(O[30]), .Z(n313) );
  ND2SVTX4 U555 ( .A(O[31]), .B(n264), .Z(n338) );
  NR2SVTX6 U556 ( .A(n237), .B(n236), .Z(n367) );
  CTIVSVTX4 U557 ( .A(O[31]), .Z(n304) );
  AO21SVTX2 U558 ( .A(N[22]), .B(n539), .C(n261), .D(n220), .Z(n240) );
  CTIVSVTX2 U559 ( .A(n261), .Z(n262) );
  IVSVTX2 U560 ( .A(N[31]), .Z(n215) );
  CTIVSVTX2 U561 ( .A(N[16]), .Z(n270) );
  CTIVSVTX2 U562 ( .A(N[1]), .Z(n330) );
  CTIVSVTX4 U563 ( .A(N[15]), .Z(n281) );
  AO7SVTX6 U564 ( .A(n793), .B(n795), .C(n794), .Z(n898) );
  B_ND2SVTX2 U565 ( .A(n794), .B(n698), .Z(n796) );
  B_ND2SVTX2 U566 ( .A(n808), .B(n807), .Z(n810) );
  B_ND2SVTX2 U567 ( .A(n798), .B(n797), .Z(n800) );
  CTIVSVTX2 U568 ( .A(n798), .Z(n787) );
  B_ND2SVTX2 U569 ( .A(n803), .B(n802), .Z(n805) );
  B_ND2SVTX2 U570 ( .A(n912), .B(n911), .Z(n913) );
  B_ND2SVTX2 U571 ( .A(n813), .B(n812), .Z(n814) );
  B_ND2SVTX2 U572 ( .A(n916), .B(n915), .Z(n918) );
  AO6SVTX2 U573 ( .A(n213), .B(n818), .C(n737), .Z(n815) );
  B_ND2SVTX2 U574 ( .A(n816), .B(n213), .Z(n817) );
  CTIVSVTX2 U575 ( .A(n816), .Z(n737) );
  B_ND2SVTX2 U576 ( .A(n897), .B(n896), .Z(n901) );
  B_ND2SVTX2 U577 ( .A(n776), .B(n775), .Z(n803) );
  FAS1SVTX2 U578 ( .A(n760), .B(n759), .CI(n758), .CO(n765), .Z(n761) );
  B_ND2SVTX1 U579 ( .A(n895), .B(n894), .Z(n897) );
  B_ND2SVTX2 U580 ( .A(n754), .B(n753), .Z(n813) );
  OR2SVTX0H U581 ( .A(n895), .B(n894), .Z(n896) );
  AO7CSVTX4 U582 ( .A(n752), .B(n777), .C(n712), .Z(n759) );
  FAS1SVTX2 U583 ( .A(n768), .B(n767), .CI(n766), .CO(n773), .Z(n764) );
  B_ND2SVTX2 U584 ( .A(n703), .B(n722), .Z(n894) );
  FAS1SVTX2 U585 ( .A(n757), .B(n756), .CI(n755), .CO(n762), .Z(n753) );
  AO6SVTX2 U586 ( .A(n750), .B(n692), .C(n711), .Z(n722) );
  AO6NSVTX2 U587 ( .A(n752), .B(n892), .C(n751), .Z(n755) );
  B_ND2SVTX2 U588 ( .A(n691), .B(n892), .Z(n703) );
  AO7SVTX6 U589 ( .A(n838), .B(n562), .C(n561), .Z(n653) );
  AO7SVTX4 U590 ( .A(n860), .B(n510), .C(n509), .Z(n843) );
  B_ND2SVTX2 U591 ( .A(n674), .B(n673), .Z(n676) );
  AO7SVTX2 U592 ( .A(n837), .B(n556), .C(n836), .Z(n560) );
  B_ND2SVTX1 U593 ( .A(n558), .B(n559), .Z(n536) );
  AO6SVTX4 U594 ( .A(n820), .B(n433), .C(n532), .Z(n837) );
  B_ND2SVTX1 U595 ( .A(n826), .B(n825), .Z(n830) );
  B_ND2SVTX1 U596 ( .A(n904), .B(n903), .Z(n906) );
  B_ND2SVTX1 U597 ( .A(n836), .B(n835), .Z(n841) );
  B_ND2SVTX1 U598 ( .A(n873), .B(n872), .Z(n875) );
  B_ND2SVTX2 U599 ( .A(n720), .B(n718), .Z(n727) );
  B_ND2SVTX2 U600 ( .A(n433), .B(n821), .Z(n839) );
  B_ND2SVTX2 U601 ( .A(n700), .B(n699), .Z(n740) );
  B_ND2SVTX1 U602 ( .A(n908), .B(n907), .Z(n910) );
  B_ND2SVTX2 U603 ( .A(n710), .B(n708), .Z(n678) );
  B_ND2SVTX1 U604 ( .A(n650), .B(n652), .Z(n563) );
  AO7SVTX2 U605 ( .A(n480), .B(n479), .C(n478), .Z(n883) );
  B_ND2SVTX1 U606 ( .A(n832), .B(n831), .Z(n834) );
  B_ND2SVTX2 U607 ( .A(n529), .B(n528), .Z(n826) );
  B_ND2SVTX2 U608 ( .A(n554), .B(n553), .Z(n650) );
  B_ND2SVTX1 U609 ( .A(n877), .B(n876), .Z(n879) );
  B_ND2SVTX1 U610 ( .A(n432), .B(n425), .Z(n558) );
  B_ND2SVTX1 U611 ( .A(n842), .B(n212), .Z(n848) );
  B_ND2SVTX1 U612 ( .A(n882), .B(n881), .Z(n885) );
  B_ND2SVTX2 U613 ( .A(n534), .B(n533), .Z(n836) );
  B_ND2SVTX2 U614 ( .A(n512), .B(n511), .Z(n873) );
  IVSVTX0H U615 ( .A(n827), .Z(n831) );
  B_ND2SVTX2 U616 ( .A(n655), .B(n654), .Z(n904) );
  B_ND2SVTX2 U617 ( .A(n858), .B(n862), .Z(n510) );
  B_ND2SVTX1 U618 ( .A(n850), .B(n849), .Z(n852) );
  B_ND2SVTX2 U619 ( .A(n531), .B(n530), .Z(n819) );
  B_ND2SVTX1 U620 ( .A(n859), .B(n858), .Z(n864) );
  CTIVSVTX2 U621 ( .A(n850), .Z(n846) );
  OR2SVTX4 U622 ( .A(n531), .B(n530), .Z(n433) );
  B_ND2SVTX1 U623 ( .A(n854), .B(n853), .Z(n857) );
  B_ND2SVTX1 U624 ( .A(n888), .B(n887), .Z(n890) );
  B_ND2SVTX2 U625 ( .A(n849), .B(n212), .Z(n523) );
  B_ND2SVTX2 U626 ( .A(n660), .B(n630), .Z(n631) );
  OR2SVTX2 U627 ( .A(n520), .B(n519), .Z(n212) );
  B_ND2SVTX2 U628 ( .A(n507), .B(n506), .Z(n859) );
  NR2SVTX2 U629 ( .A(n527), .B(n526), .Z(n827) );
  B_ND2SVTX2 U630 ( .A(n527), .B(n526), .Z(n832) );
  B_ND2SVTX2 U631 ( .A(n514), .B(n513), .Z(n854) );
  AO7SVTX2 U632 ( .A(n888), .B(n880), .C(n882), .Z(n489) );
  B_ND2SVTX2 U633 ( .A(n518), .B(n517), .Z(n850) );
  B_ND2SVTX2 U634 ( .A(n660), .B(n634), .Z(n635) );
  B_ND2SVTX2 U635 ( .A(n660), .B(n637), .Z(n638) );
  B_ND2SVTX2 U636 ( .A(n520), .B(n519), .Z(n842) );
  B_ND2SVTX2 U637 ( .A(n503), .B(n502), .Z(n877) );
  B_ND2SVTX2 U638 ( .A(n505), .B(n504), .Z(n867) );
  B_ND2SVTX2 U639 ( .A(n661), .B(n660), .Z(n662) );
  B_ND2SVTX2 U640 ( .A(n488), .B(n487), .Z(n882) );
  B_ND2SVTX2 U641 ( .A(n463), .B(n462), .Z(n469) );
  B_ND2SVTX2 U642 ( .A(n486), .B(n485), .Z(n888) );
  F_EOSVTX2 U643 ( .A(n432), .B(n431), .Z(n437) );
  B_ND2SVTX2 U644 ( .A(n656), .B(n660), .Z(n657) );
  F_ENSVTX2 U645 ( .A(n554), .B(n660), .Z(n443) );
  B_ND2SVTX1 U646 ( .A(n550), .B(n660), .Z(n551) );
  B_ND2SVTX2 U647 ( .A(n491), .B(n435), .Z(n436) );
  B_ND2SVTX2 U648 ( .A(n491), .B(n439), .Z(n440) );
  B_ND2SVTX2 U649 ( .A(n445), .B(n491), .Z(n446) );
  B_ND2SVTX2 U650 ( .A(n455), .B(n491), .Z(n456) );
  B_ND2SVTX2 U651 ( .A(n447), .B(n491), .Z(n448) );
  ENSVTX0H U652 ( .A(n507), .B(n483), .Z(n499) );
  BFSVTX6 U653 ( .A(n683), .Z(n691) );
  B_ND2SVTX2 U654 ( .A(n445), .B(n407), .Z(n408) );
  B_ND2SVTX2 U655 ( .A(n626), .B(n640), .Z(n627) );
  IVSVTX4 U656 ( .A(n893), .Z(n683) );
  B_ND2SVTX2 U657 ( .A(n588), .B(n587), .Z(n589) );
  B_ND2SVTX2 U658 ( .A(n586), .B(n585), .Z(n636) );
  NR2SVTX2 U659 ( .A(n752), .B(n692), .Z(n751) );
  CTIVSVTX2 U660 ( .A(n655), .Z(n421) );
  B_ND2SVTX2 U661 ( .A(n360), .B(n359), .Z(n493) );
  B_ND2SVTX2 U662 ( .A(n391), .B(n428), .Z(n406) );
  F_IVSVTX1 U663 ( .A(n531), .Z(n404) );
  AO7SVTX4 U664 ( .A(n272), .B(n573), .C(n567), .Z(n697) );
  F_IVSVTX1 U665 ( .A(n503), .Z(n359) );
  F_IVSVTX1 U666 ( .A(n488), .Z(n470) );
  AO2ASVTX2 U667 ( .C(n415), .D(n392), .A(n321), .B(n583), .Z(n322) );
  AO39SVTX2 U668 ( .A(n599), .B(n591), .C(n600), .D(n570), .E(n569), .F(n568), 
        .Z(n582) );
  F_IVSVTX1 U669 ( .A(n505), .Z(n360) );
  CTIVSVTX2 U670 ( .A(n518), .Z(n369) );
  AO1SVTX2 U671 ( .A(n278), .B(n385), .C(n269), .D(n268), .Z(n323) );
  MUX21NSVTX2 U672 ( .A(n352), .B(n351), .S(O[28]), .Z(n505) );
  CTIVSVTX2 U673 ( .A(n604), .Z(n412) );
  CTIVSVTX2 U674 ( .A(n621), .Z(n592) );
  CTIVSVTX2 U675 ( .A(n591), .Z(n611) );
  AO2SVTX2 U676 ( .A(N[6]), .B(n366), .C(n393), .D(O[29]), .Z(n373) );
  AO6ABSVTX2 U677 ( .A(n283), .B(n542), .C(n277), .Z(n616) );
  MUX21NSVTX2 U678 ( .A(N[2]), .B(N[3]), .S(O[27]), .Z(n331) );
  AO6ABSVTX2 U679 ( .A(n275), .B(n542), .C(n274), .Z(n621) );
  AO2SVTX2 U680 ( .A(N[7]), .B(n366), .C(n385), .D(O[29]), .Z(n375) );
  B_ND2SVTX2 U681 ( .A(N[0]), .B(n313), .Z(n295) );
  ND4ABSVTX6 U682 ( .A(n240), .B(n239), .C(n238), .D(n367), .Z(n272) );
  B_ND2SVTX2 U683 ( .A(n270), .B(n306), .Z(n226) );
  NR4SVTX4 U684 ( .A(N[23]), .B(N[21]), .C(N[22]), .D(N[20]), .Z(n245) );
  CTIVSVTX2 U685 ( .A(N[6]), .Z(n345) );
  IVSVTX0H U686 ( .A(N[0]), .Z(n329) );
  CTIVSVTX2 U687 ( .A(N[7]), .Z(n343) );
  CTIVSVTX2 U688 ( .A(N[22]), .Z(n308) );
  CTIVSVTX2 U689 ( .A(N[5]), .Z(n538) );
  NR2SVTX2 U690 ( .A(n432), .B(n425), .Z(n557) );
  AO11NSVTX4 U691 ( .A(n655), .B(n684), .C(n683), .D(n442), .E(n444), .F(n552), 
        .Z(n425) );
  AO11NSVTX2 U692 ( .A(n477), .B(n704), .C(n691), .D(n464), .E(n701), .F(n210), 
        .Z(n465) );
  IVSVTX4 U693 ( .A(n265), .Z(O[30]) );
  NR2SVTX2 U694 ( .A(n721), .B(n711), .Z(n712) );
  NR2SVTX2 U695 ( .A(n376), .B(n375), .Z(n377) );
  AO3SVTX2 U696 ( .A(n743), .B(n784), .C(n722), .D(n721), .Z(n767) );
  F_ENSVTX2 U697 ( .A(n514), .B(n491), .Z(n500) );
  AO11NSVTX4 U698 ( .A(n710), .B(n684), .C(n683), .D(n665), .E(n444), .F(n664), 
        .Z(n747) );
  EOSVTX4 U699 ( .A(n901), .B(n900), .Z(O[26]) );
  ND2SVTX4 U700 ( .A(n697), .B(n689), .Z(n731) );
  ND2SVTX4 U701 ( .A(n899), .B(n898), .Z(n900) );
  ENSVTX4 U702 ( .A(n690), .B(n689), .Z(n750) );
  NR2SVTX2 U703 ( .A(n824), .B(n827), .Z(n821) );
  AO7SVTX2 U704 ( .A(n844), .B(n523), .C(n522), .Z(n524) );
  AO11NSVTX1 U705 ( .A(n514), .B(n704), .C(n691), .D(n500), .E(n701), .F(n492), 
        .Z(n506) );
  AO11NSVTX2 U706 ( .A(n534), .B(n704), .C(n691), .D(n441), .E(n444), .F(n437), 
        .Z(n528) );
  AO4SVTX1 U707 ( .A(n540), .B(n306), .C(n344), .D(n537), .Z(n274) );
  CTIVSVTX2 U708 ( .A(n375), .Z(n372) );
  AO11NSVTX1 U709 ( .A(n503), .B(n704), .C(n691), .D(n482), .E(n701), .F(n484), 
        .Z(n485) );
  AO11NSVTX2 U710 ( .A(n512), .B(n704), .C(n691), .D(n501), .E(n701), .F(n500), 
        .Z(n504) );
  AO11NSVTX1 U711 ( .A(n554), .B(n684), .C(n683), .D(n443), .E(n444), .F(n442), 
        .Z(n533) );
  AO7SVTX4 U712 ( .A(n417), .B(n323), .C(n273), .Z(n432) );
  CTIVSVTX2 U713 ( .A(n819), .Z(n532) );
  F_MUX21NSVTX1 U714 ( .A(n330), .B(n344), .S(n583), .Z(n332) );
  AO11NSVTX1 U715 ( .A(n488), .B(n704), .C(n691), .D(n470), .E(n701), .F(n482), 
        .Z(n476) );
  F_ND2SVTX0H U716 ( .A(n714), .B(n713), .Z(n716) );
  AO6SVTX1 U717 ( .A(n212), .B(n846), .C(n521), .Z(n522) );
  CTIVSVTX4 U718 ( .A(N[14]), .Z(n310) );
  AO7ASVTX4 U719 ( .A(n263), .B(O[31]), .C(n262), .Z(n264) );
  CTIVSVTX4 U720 ( .A(N[18]), .Z(n306) );
  EOSVTX0H U721 ( .A(n890), .B(n889), .Z(O[0]) );
  ENSVTX0H U722 ( .A(n885), .B(n884), .Z(O[1]) );
  ENSVTX0H U723 ( .A(n879), .B(n878), .Z(O[2]) );
  EOSVTX0H U724 ( .A(n871), .B(n870), .Z(O[3]) );
  EOSVTX0H U725 ( .A(n864), .B(n863), .Z(O[4]) );
  EOSVTX0H U726 ( .A(n875), .B(n874), .Z(O[5]) );
  ENSVTX0H U727 ( .A(n857), .B(n856), .Z(O[6]) );
  ENSVTX0H U728 ( .A(n852), .B(n851), .Z(O[7]) );
  EOSVTX0H U729 ( .A(n848), .B(n847), .Z(O[8]) );
  ENSVTX0H U730 ( .A(n834), .B(n833), .Z(O[9]) );
  EOSVTX0H U731 ( .A(n830), .B(n829), .Z(O[10]) );
  EOSVTX0H U732 ( .A(n823), .B(n822), .Z(O[11]) );
  ENSVTX0H U733 ( .A(n841), .B(n840), .Z(O[12]) );
  EOSVTX0H U734 ( .A(n536), .B(n535), .Z(O[13]) );
  ENSVTX0H U735 ( .A(n910), .B(n909), .Z(O[16]) );
  OR2SVTX2 U736 ( .A(n735), .B(n734), .Z(n213) );
  F_IVSVTX0H U737 ( .A(n264), .Z(n265) );
  ND2SVTX4 U738 ( .A(n298), .B(n215), .Z(n216) );
  NR3SVTX8 U739 ( .A(N[30]), .B(N[29]), .C(n216), .Z(n346) );
  IVSVTX0H U740 ( .A(N[26]), .Z(n219) );
  IVSVTX0H U741 ( .A(N[29]), .Z(n287) );
  AO8SVTX1 U742 ( .A(N[25]), .B(n219), .C(n346), .D(n218), .Z(n220) );
  NR2ASVTX6 U743 ( .A(n245), .B(n261), .Z(n229) );
  NR3ABSVTX2 U744 ( .A(N[17]), .B(n306), .C(n250), .Z(n239) );
  NR4SVTX2 U745 ( .A(N[4]), .B(N[5]), .C(N[6]), .D(N[7]), .Z(n241) );
  NR2SVTX2 U746 ( .A(N[11]), .B(N[9]), .Z(n223) );
  NR2SVTX2 U747 ( .A(N[8]), .B(N[10]), .Z(n222) );
  NR2SVTX2 U748 ( .A(N[13]), .B(N[12]), .Z(n221) );
  ND3SVTX4 U749 ( .A(n281), .B(n310), .C(n221), .Z(n242) );
  NR3SVTX2 U750 ( .A(N[2]), .B(n330), .C(n251), .Z(n228) );
  IVSVTX2 U751 ( .A(n242), .Z(n252) );
  ND4ABCSVTX8 U752 ( .A(N[17]), .B(N[19]), .C(n226), .D(n229), .Z(O[31]) );
  AO7SVTX2 U753 ( .A(n228), .B(n227), .C(n304), .Z(n238) );
  F_AN2SVTX2 U754 ( .A(N[19]), .B(n229), .Z(n232) );
  NR2ASVTX1 U755 ( .A(N[23]), .B(n261), .Z(n230) );
  AO1SVTX2 U756 ( .A(n346), .B(N[27]), .C(N[31]), .D(n230), .Z(n231) );
  F_ND2ASVTX2 U757 ( .A(n232), .B(n231), .Z(n237) );
  AO6SVTX1 U758 ( .A(n252), .B(N[11]), .C(N[15]), .Z(n233) );
  AO7SVTX2 U759 ( .A(n343), .B(n263), .C(n233), .Z(n235) );
  NR2ASVTX2 U760 ( .A(N[3]), .B(n251), .Z(n234) );
  AO6ABSVTX2 U761 ( .A(n235), .B(n234), .C(O[31]), .Z(n236) );
  IVSVTX0H U762 ( .A(n241), .Z(n243) );
  NR2SVTX2 U763 ( .A(n245), .B(n261), .Z(n246) );
  AO6SVTX1 U764 ( .A(n346), .B(N[26]), .C(N[30]), .Z(n249) );
  NR2ASVTX2 U765 ( .A(N[18]), .B(n250), .Z(n259) );
  AO6SVTX1 U766 ( .A(n252), .B(N[10]), .C(N[14]), .Z(n253) );
  AO7SVTX2 U767 ( .A(n345), .B(n263), .C(n253), .Z(n254) );
  AO6SVTX2 U768 ( .A(N[2]), .B(n255), .C(n254), .Z(n256) );
  F_ND2ASVTX2 U769 ( .A(n256), .B(n304), .Z(n257) );
  ND4ABCSVTX8 U770 ( .A(n260), .B(n259), .C(n258), .D(n367), .Z(O[28]) );
  OR2SVTX4 U771 ( .A(n304), .B(n264), .Z(n542) );
  IVSVTX0H U772 ( .A(N[9]), .Z(n337) );
  IVSVTX0H U773 ( .A(N[17]), .Z(n266) );
  AO6ABSVTX2 U774 ( .A(n337), .B(n542), .C(n267), .Z(n620) );
  AO4SVTX1 U775 ( .A(n620), .B(n569), .C(n599), .D(n370), .Z(n268) );
  IVSVTX0H U776 ( .A(N[12]), .Z(n300) );
  AO4SVTX1 U777 ( .A(n542), .B(n345), .C(n310), .D(n540), .Z(n414) );
  IVSVTX0H U778 ( .A(N[8]), .Z(n339) );
  AO4SVTX1 U779 ( .A(n540), .B(n270), .C(n329), .D(n537), .Z(n271) );
  AO6ABSVTX2 U780 ( .A(n339), .B(n542), .C(n271), .Z(n604) );
  AO39SVTX2 U781 ( .A(n599), .B(n320), .C(n600), .D(n546), .E(n569), .F(n604), 
        .Z(n389) );
  AO2SVTX2 U782 ( .A(n389), .B(n420), .C(n211), .D(n393), .Z(n273) );
  IVSVTX4 U783 ( .A(n599), .Z(n612) );
  IVSVTX4 U784 ( .A(n600), .Z(n610) );
  IVSVTX0H U785 ( .A(N[19]), .Z(n276) );
  AO4SVTX1 U786 ( .A(n214), .B(n370), .C(n320), .D(n397), .Z(n279) );
  AO6SVTX1 U787 ( .A(n419), .B(n583), .C(n279), .Z(n280) );
  IVSVTX2 U788 ( .A(n313), .Z(n301) );
  NR2ASVTX1 U789 ( .A(N[19]), .B(O[30]), .Z(n282) );
  AO1ABSVTX1 U790 ( .A(O[31]), .B(n283), .C(N[27]), .D(n282), .Z(n284) );
  AO20SVTX2 U791 ( .A(n342), .B(n301), .C(n284), .D(n341), .Z(n286) );
  NR2ASVTX1 U792 ( .A(N[23]), .B(n363), .Z(n285) );
  AO1SVTX2 U793 ( .A(n341), .B(n597), .C(n286), .D(n285), .Z(n564) );
  IVSVTX2 U794 ( .A(n537), .Z(n410) );
  AO7SVTX1 U795 ( .A(n539), .B(O[30]), .C(n287), .Z(n288) );
  AO6SVTX1 U796 ( .A(n410), .B(N[13]), .C(n288), .Z(n289) );
  AO7SVTX1 U797 ( .A(n538), .B(n301), .C(n289), .Z(n292) );
  NR2ASVTX1 U798 ( .A(N[17]), .B(O[30]), .Z(n290) );
  AO1ABSVTX1 U799 ( .A(O[31]), .B(n337), .C(N[25]), .D(n290), .Z(n291) );
  AO2SVTX2 U800 ( .A(n614), .B(n292), .C(n612), .D(n574), .Z(n293) );
  AO7SVTX2 U801 ( .A(O[28]), .B(n564), .C(n293), .Z(n319) );
  IVSVTX0H U802 ( .A(N[24]), .Z(n294) );
  AO7SVTX1 U803 ( .A(n339), .B(O[31]), .C(n294), .Z(n297) );
  NR2ASVTX1 U804 ( .A(N[16]), .B(O[30]), .Z(n296) );
  ND3ABSVTX2 U805 ( .A(n297), .B(n296), .C(n295), .Z(n615) );
  IVSVTX0H U806 ( .A(N[20]), .Z(n299) );
  AO7SVTX1 U807 ( .A(n299), .B(n542), .C(n298), .Z(n303) );
  IVSVTX0H U808 ( .A(N[4]), .Z(n340) );
  AO4SVTX1 U809 ( .A(n301), .B(n340), .C(n537), .D(n300), .Z(n302) );
  AO1SVTX2 U810 ( .A(n341), .B(n615), .C(n303), .D(n302), .Z(n317) );
  AO6SVTX1 U811 ( .A(n304), .B(N[10]), .C(N[26]), .Z(n305) );
  AO7SVTX1 U812 ( .A(n306), .B(O[30]), .C(n305), .Z(n307) );
  AO6ASVTX2 U813 ( .A(n344), .B(n313), .C(n307), .Z(n568) );
  AO4SVTX2 U814 ( .A(n317), .B(n379), .C(n568), .D(n600), .Z(n566) );
  AO4SVTX1 U815 ( .A(n540), .B(n308), .C(n345), .D(n537), .Z(n309) );
  AO2ABSVTX2 U816 ( .C(n417), .D(n566), .A(n591), .B(n397), .Z(n311) );
  ND2SVTX4 U817 ( .A(n312), .B(n311), .Z(n632) );
  F_AO2SVTX1 U818 ( .A(n411), .B(N[22]), .C(N[6]), .D(n313), .Z(n315) );
  AO6SVTX1 U819 ( .A(n410), .B(N[14]), .C(N[30]), .Z(n314) );
  AO3SVTX1 U820 ( .A(n568), .B(n599), .C(n315), .D(n314), .Z(n316) );
  NR2SVTX2 U821 ( .A(n325), .B(n324), .Z(n466) );
  NR2SVTX2 U822 ( .A(n466), .B(n463), .Z(n328) );
  NR2ASVTX2 U823 ( .A(n209), .B(n600), .Z(n354) );
  IVSVTX2 U824 ( .A(n354), .Z(n576) );
  NR2SVTX2 U825 ( .A(n477), .B(n472), .Z(n327) );
  AO4SVTX1 U826 ( .A(n346), .B(n340), .C(n329), .D(n363), .Z(n356) );
  AO4SVTX1 U827 ( .A(n346), .B(n538), .C(n330), .D(n363), .Z(n349) );
  IVSVTX0H U828 ( .A(n356), .Z(n334) );
  NR2ASVTX1 U829 ( .A(N[3]), .B(n272), .Z(n353) );
  F_AO2SVTX1 U830 ( .A(n354), .B(n332), .C(n598), .D(n353), .Z(n333) );
  AO7SVTX2 U831 ( .A(n334), .B(n367), .C(n333), .Z(n486) );
  NR2SVTX2 U832 ( .A(n336), .B(n335), .Z(n460) );
  AO4SVTX2 U833 ( .A(n399), .B(n341), .C(n538), .D(n363), .Z(n378) );
  AO4SVTX2 U834 ( .A(n398), .B(n341), .C(n340), .D(n363), .Z(n348) );
  MUX21NSVTX2 U835 ( .A(n378), .B(n348), .S(n417), .Z(n368) );
  AO4SVTX1 U836 ( .A(n346), .B(n343), .C(n342), .D(n363), .Z(n347) );
  AO4SVTX1 U837 ( .A(n346), .B(n345), .C(n344), .D(n363), .Z(n350) );
  MUX21NSVTX2 U838 ( .A(n347), .B(n350), .S(n417), .Z(n351) );
  MUX21NSVTX2 U839 ( .A(n348), .B(n347), .S(n417), .Z(n365) );
  MUX21NSVTX2 U840 ( .A(n350), .B(n349), .S(n417), .Z(n358) );
  F_AN2SVTX2 U841 ( .A(n379), .B(n583), .Z(n355) );
  F_AO2SVTX1 U842 ( .A(n356), .B(n355), .C(n354), .D(n353), .Z(n357) );
  AO7SVTX4 U843 ( .A(n379), .B(n358), .C(n357), .Z(n503) );
  NR3ABSVTX2 U844 ( .A(n361), .B(n495), .C(n493), .Z(n362) );
  ND2SVTX4 U845 ( .A(n460), .B(n362), .Z(n426) );
  IVSVTX0H U846 ( .A(n378), .Z(n364) );
  AO39SVTX2 U847 ( .A(n365), .B(O[28]), .C(n376), .D(n364), .E(n367), .F(n373), 
        .Z(n514) );
  AO39SVTX2 U848 ( .A(n368), .B(O[28]), .C(n367), .D(n375), .E(n376), .F(n373), 
        .Z(n518) );
  AO11SVTX2 U849 ( .A(n372), .B(n379), .C(n413), .D(n614), .E(n371), .F(n612), 
        .Z(n396) );
  AO11SVTX2 U850 ( .A(n374), .B(n379), .C(n392), .D(n614), .E(n394), .F(n612), 
        .Z(n381) );
  MUX21NSVTX2 U851 ( .A(n396), .B(n381), .S(n420), .Z(n527) );
  AO8SVTX1 U852 ( .A(n379), .B(n420), .C(n378), .D(n377), .Z(n380) );
  NR2SVTX2 U853 ( .A(n451), .B(n384), .Z(n445) );
  AO11SVTX4 U854 ( .A(n386), .B(n614), .C(n385), .D(n612), .E(n413), .F(n610), 
        .Z(n401) );
  IVSVTX0H U855 ( .A(n393), .Z(n387) );
  AO4SVTX1 U856 ( .A(n214), .B(n387), .C(n399), .D(n397), .Z(n388) );
  AO6SVTX2 U857 ( .A(n389), .B(n583), .C(n388), .Z(n390) );
  AO11SVTX2 U858 ( .A(n414), .B(n614), .C(n393), .D(n612), .E(n392), .F(n610), 
        .Z(n403) );
  AO2ASVTX4 U859 ( .C(n415), .D(n394), .A(n403), .B(O[27]), .Z(n395) );
  AO4SVTX1 U860 ( .A(n214), .B(n399), .C(n398), .D(n397), .Z(n400) );
  AO6ABSVTX2 U861 ( .A(n417), .B(n401), .C(n400), .Z(n402) );
  AO7SVTX4 U862 ( .A(n403), .B(O[27]), .C(n402), .Z(n531) );
  NR2SVTX2 U863 ( .A(n406), .B(n434), .Z(n407) );
  ND2SVTX4 U864 ( .A(n422), .B(n660), .Z(n409) );
  F_EOSVTX2 U865 ( .A(n655), .B(n409), .Z(n442) );
  F_AO2SVTX1 U866 ( .A(n415), .B(n414), .C(n211), .D(n413), .Z(n416) );
  F_EOSVTX2 U867 ( .A(n670), .B(n424), .Z(n552) );
  IVSVTX2 U868 ( .A(n445), .Z(n438) );
  F_IVSVTX0H U869 ( .A(n434), .Z(n427) );
  ND2SVTX2 U870 ( .A(n428), .B(n427), .Z(n429) );
  NR2SVTX2 U871 ( .A(n438), .B(n429), .Z(n430) );
  ND2SVTX2 U872 ( .A(n491), .B(n430), .Z(n431) );
  NR2SVTX2 U873 ( .A(n434), .B(n438), .Z(n435) );
  F_EOSVTX2 U874 ( .A(n534), .B(n436), .Z(n441) );
  NR2SVTX2 U875 ( .A(n529), .B(n528), .Z(n824) );
  NR2SVTX2 U876 ( .A(n529), .B(n438), .Z(n439) );
  AO11NSVTX4 U877 ( .A(n531), .B(n704), .C(n691), .D(n449), .E(n701), .F(n441), 
        .Z(n526) );
  NR2SVTX2 U878 ( .A(n534), .B(n533), .Z(n556) );
  IVSVTX0H U879 ( .A(n556), .Z(n835) );
  NR2SVTX0H U880 ( .A(n520), .B(n451), .Z(n447) );
  AO11NSVTX2 U881 ( .A(n701), .B(n450), .C(n684), .D(n527), .E(n691), .F(n454), 
        .Z(n517) );
  OR2SVTX2 U882 ( .A(n518), .B(n517), .Z(n849) );
  AO11NSVTX4 U883 ( .A(n529), .B(n704), .C(n691), .D(n450), .E(n701), .F(n449), 
        .Z(n519) );
  IVSVTX0H U884 ( .A(n451), .Z(n452) );
  AO11NSVTX4 U885 ( .A(n520), .B(n704), .C(n691), .D(n457), .E(n701), .F(n454), 
        .Z(n513) );
  OR2SVTX2 U886 ( .A(n514), .B(n513), .Z(n853) );
  F_EOSVTX2 U887 ( .A(n518), .B(n456), .Z(n492) );
  F_AO2SVTX1 U888 ( .A(n457), .B(n701), .C(n704), .D(n518), .Z(n458) );
  NR2SVTX2 U889 ( .A(n512), .B(n511), .Z(n855) );
  NR2SVTX2 U890 ( .A(n523), .B(n845), .Z(n525) );
  IVSVTX2 U891 ( .A(n460), .Z(n497) );
  EOSVTX0H U892 ( .A(n503), .B(n497), .Z(n482) );
  NR2SVTX2 U893 ( .A(n477), .B(n476), .Z(n480) );
  IVSVTX0H U894 ( .A(n472), .Z(n461) );
  IVSVTX0H U895 ( .A(n477), .Z(n464) );
  AO11NSVTX1 U896 ( .A(n472), .B(n704), .C(n691), .D(n461), .E(n701), .F(n464), 
        .Z(n462) );
  NR2SVTX2 U897 ( .A(n466), .B(n465), .Z(n468) );
  B_ND2SVTX1 U898 ( .A(n466), .B(n465), .Z(n467) );
  AO7SVTX2 U899 ( .A(n469), .B(n468), .C(n467), .Z(n475) );
  AO11NSVTX1 U900 ( .A(n486), .B(n704), .C(n691), .D(n210), .E(n701), .F(n470), 
        .Z(n471) );
  OR2SVTX2 U901 ( .A(n472), .B(n471), .Z(n474) );
  F_AN2SVTX2 U902 ( .A(n472), .B(n471), .Z(n473) );
  AO6SVTX2 U903 ( .A(n475), .B(n474), .C(n473), .Z(n479) );
  NR2SVTX2 U904 ( .A(n503), .B(n497), .Z(n481) );
  ENSVTX0H U905 ( .A(n505), .B(n481), .Z(n484) );
  NR2SVTX2 U906 ( .A(n486), .B(n485), .Z(n886) );
  NR2SVTX2 U907 ( .A(n493), .B(n497), .Z(n483) );
  AO11NSVTX2 U908 ( .A(n505), .B(n704), .C(n691), .D(n484), .E(n701), .F(n499), 
        .Z(n487) );
  NR2SVTX2 U909 ( .A(n488), .B(n487), .Z(n880) );
  NR2SVTX2 U910 ( .A(n886), .B(n880), .Z(n490) );
  OR2SVTX2 U911 ( .A(n507), .B(n506), .Z(n858) );
  IVSVTX0H U912 ( .A(n493), .Z(n494) );
  NR2SVTX2 U913 ( .A(n497), .B(n496), .Z(n498) );
  NR2SVTX2 U914 ( .A(n503), .B(n502), .Z(n868) );
  NR2SVTX2 U915 ( .A(n505), .B(n504), .Z(n865) );
  NR2SVTX2 U916 ( .A(n868), .B(n865), .Z(n862) );
  AO7SVTX2 U917 ( .A(n877), .B(n865), .C(n867), .Z(n861) );
  AO6SVTX2 U918 ( .A(n861), .B(n858), .C(n508), .Z(n509) );
  F_IVSVTX0H U919 ( .A(n854), .Z(n515) );
  AO6SVTX1 U920 ( .A(n853), .B(n516), .C(n515), .Z(n844) );
  AO7SVTX4 U921 ( .A(n832), .B(n824), .C(n826), .Z(n820) );
  AO8SVTX1 U922 ( .A(n555), .B(n835), .C(n833), .D(n560), .Z(n535) );
  AO4SVTX1 U923 ( .A(n540), .B(n539), .C(n538), .D(n537), .Z(n541) );
  IVSVTX0H U924 ( .A(n620), .Z(n545) );
  AO11SVTX2 U925 ( .A(n579), .B(n614), .C(n545), .D(n612), .E(n544), .F(n610), 
        .Z(n596) );
  AO4SVTX1 U926 ( .A(n214), .B(n593), .C(n546), .D(n397), .Z(n547) );
  AO6ABSVTX1 U927 ( .A(n417), .B(n596), .C(n547), .Z(n548) );
  AO7SVTX2 U928 ( .A(n549), .B(n272), .C(n548), .Z(n749) );
  NR2SVTX0H U929 ( .A(n670), .B(n590), .Z(n550) );
  AO11NSVTX2 U930 ( .A(n670), .B(n684), .C(n683), .D(n552), .E(n444), .F(n649), 
        .Z(n553) );
  OR2SVTX2 U931 ( .A(n554), .B(n553), .Z(n652) );
  ND3ABSVTX2 U932 ( .A(n557), .B(n556), .C(n555), .Z(n562) );
  AO6CSVTX2 U933 ( .A(n560), .B(n559), .C(n558), .Z(n561) );
  ENSVTX0H U934 ( .A(n563), .B(n653), .Z(O[14]) );
  AO4SVTX1 U935 ( .A(n214), .B(n591), .C(n601), .D(n397), .Z(n565) );
  IVSVTX0H U936 ( .A(n615), .Z(n570) );
  AO4SVTX1 U937 ( .A(n580), .B(n397), .C(n601), .D(n214), .Z(n571) );
  AO6SVTX1 U938 ( .A(n417), .B(n582), .C(n571), .Z(n572) );
  IVSVTX0H U939 ( .A(N[23]), .Z(n577) );
  AO7SVTX1 U940 ( .A(n577), .B(n576), .C(n575), .Z(n578) );
  AO4SVTX1 U941 ( .A(n580), .B(n214), .C(n616), .D(n397), .Z(n581) );
  AO4SVTX1 U942 ( .A(n214), .B(n604), .C(n593), .D(n397), .Z(n594) );
  AO6ABSVTX1 U943 ( .A(n420), .B(n607), .C(n594), .Z(n595) );
  AO7SVTX2 U944 ( .A(n596), .B(O[27]), .C(n595), .Z(n746) );
  F_AO2SVTX1 U945 ( .A(n598), .B(N[23]), .C(n614), .D(n597), .Z(n603) );
  AO4SVTX1 U946 ( .A(n601), .B(n600), .C(n599), .D(n616), .Z(n602) );
  AO4SVTX1 U947 ( .A(n214), .B(n620), .C(n604), .D(n397), .Z(n605) );
  AO6ABSVTX1 U948 ( .A(n417), .B(n625), .C(n605), .Z(n606) );
  AO4SVTX1 U949 ( .A(n214), .B(n616), .C(n621), .D(n397), .Z(n617) );
  AO4SVTX1 U950 ( .A(n214), .B(n621), .C(n620), .D(n397), .Z(n622) );
  AO7SVTX2 U951 ( .A(n625), .B(n583), .C(n624), .Z(n720) );
  NR2SVTX2 U952 ( .A(n658), .B(n627), .Z(n628) );
  NR2SVTX2 U953 ( .A(n629), .B(n644), .Z(n630) );
  NR2SVTX2 U954 ( .A(n707), .B(n644), .Z(n634) );
  NR2SVTX2 U955 ( .A(n636), .B(n644), .Z(n637) );
  NR2SVTX2 U956 ( .A(n659), .B(n641), .Z(n642) );
  F_EOSVTX2 U957 ( .A(n700), .B(n643), .Z(n663) );
  NR2SVTX2 U958 ( .A(n710), .B(n708), .Z(n680) );
  AO11NSVTX2 U959 ( .A(n749), .B(n684), .C(n683), .D(n649), .E(n444), .F(n666), 
        .Z(n654) );
  NR2SVTX2 U960 ( .A(n655), .B(n654), .Z(n902) );
  AO6SVTX8 U961 ( .A(n653), .B(n652), .C(n651), .Z(n905) );
  AO7SVTX8 U962 ( .A(n902), .B(n905), .C(n904), .Z(n909) );
  NR2SVTX2 U963 ( .A(n746), .B(n659), .Z(n656) );
  F_EOSVTX2 U964 ( .A(n710), .B(n657), .Z(n665) );
  NR2SVTX2 U965 ( .A(n659), .B(n658), .Z(n661) );
  F_EOSVTX2 U966 ( .A(n720), .B(n662), .Z(n664) );
  NR2SVTX2 U967 ( .A(n749), .B(n747), .Z(n672) );
  AO11NSVTX4 U968 ( .A(n720), .B(n684), .C(n683), .D(n664), .E(n444), .F(n663), 
        .Z(n745) );
  NR2SVTX2 U969 ( .A(n746), .B(n745), .Z(n668) );
  AO11NSVTX4 U970 ( .A(n746), .B(n684), .C(n683), .D(n666), .E(n444), .F(n665), 
        .Z(n669) );
  OR2SVTX2 U971 ( .A(n670), .B(n669), .Z(n907) );
  NR3SVTX2 U972 ( .A(n672), .B(n668), .C(n667), .Z(n677) );
  AO1CDSVTX8 U973 ( .A(n909), .B(n677), .C(n676), .D(n675), .Z(n679) );
  AO7SVTX8 U974 ( .A(n680), .B(n679), .C(n678), .Z(n728) );
  OR2SVTX2 U975 ( .A(n720), .B(n718), .Z(n726) );
  AO6SVTX8 U976 ( .A(n728), .B(n726), .C(n685), .Z(n741) );
  AO7SVTX8 U977 ( .A(n738), .B(n741), .C(n740), .Z(n715) );
  AO11NSVTX4 U978 ( .A(n697), .B(n704), .C(n691), .D(n687), .E(n701), .F(n686), 
        .Z(n705) );
  OR2SVTX2 U979 ( .A(n694), .B(n693), .Z(n899) );
  AO3SVTX2 U980 ( .A(n731), .B(n704), .C(n703), .D(n702), .Z(n770) );
  NR2SVTX2 U981 ( .A(n776), .B(n775), .Z(n801) );
  ENSVTX0H U982 ( .A(n716), .B(n715), .Z(n717) );
  NR2ASVTX2 U983 ( .A(n717), .B(n743), .Z(n758) );
  NR2SVTX2 U984 ( .A(n765), .B(n764), .Z(n806) );
  ENSVTX0H U985 ( .A(n729), .B(n728), .Z(n730) );
  NR2ASVTX2 U986 ( .A(n730), .B(n743), .Z(n735) );
  AO7ABSVTX2 U987 ( .A(n909), .B(n907), .C(n908), .Z(n748) );
  IVSVTX0H U988 ( .A(n752), .Z(n733) );
  ND3SVTX1 U989 ( .A(n731), .B(n743), .C(n733), .Z(n732) );
  AO7SVTX2 U990 ( .A(n743), .B(n733), .C(n732), .Z(n818) );
  IVSVTX0H U991 ( .A(n734), .Z(n736) );
  F_ND2ASVTX2 U992 ( .A(n736), .B(n735), .Z(n816) );
  IVSVTX0H U993 ( .A(n738), .Z(n739) );
  EOSVTX0H U994 ( .A(n742), .B(n741), .Z(n744) );
  HA1SVTX1 U995 ( .A(n746), .B(n745), .CO(n709), .S(n757) );
  NR2SVTX2 U996 ( .A(n754), .B(n753), .Z(n811) );
  AO7SVTX4 U997 ( .A(n815), .B(n811), .C(n813), .Z(n914) );
  OR2SVTX4 U999 ( .A(n786), .B(n785), .Z(n797) );
  AO6SVTX8 U1000 ( .A(n799), .B(n797), .C(n787), .Z(n795) );
  F_ENSVTX2 U1001 ( .A(n792), .B(n898), .Z(O[25]) );
  F_EOSVTX2 U1002 ( .A(n796), .B(n795), .Z(O[24]) );
  F_EOSVTX2 U1003 ( .A(n805), .B(n804), .Z(O[22]) );
  AO6SVTX1 U1004 ( .A(n833), .B(n821), .C(n820), .Z(n822) );
  IVSVTX0H U1005 ( .A(n824), .Z(n825) );
  IVSVTX0H U1006 ( .A(n832), .Z(n828) );
  AO6SVTX1 U1007 ( .A(n833), .B(n831), .C(n828), .Z(n829) );
  AO7SVTX1 U1008 ( .A(n839), .B(n838), .C(n837), .Z(n840) );
  AO7SVTX1 U1009 ( .A(n845), .B(n874), .C(n844), .Z(n851) );
  AO6SVTX1 U1010 ( .A(n851), .B(n849), .C(n846), .Z(n847) );
  AO7SVTX1 U1011 ( .A(n855), .B(n874), .C(n873), .Z(n856) );
  AO6SVTX1 U1012 ( .A(n878), .B(n862), .C(n861), .Z(n863) );
  IVSVTX0H U1013 ( .A(n865), .Z(n866) );
  IVSVTX0H U1014 ( .A(n868), .Z(n876) );
  IVSVTX0H U1015 ( .A(n877), .Z(n869) );
  AO6SVTX1 U1016 ( .A(n878), .B(n876), .C(n869), .Z(n870) );
  IVSVTX0H U1017 ( .A(n880), .Z(n881) );
  AO7SVTX1 U1018 ( .A(n886), .B(n889), .C(n888), .Z(n884) );
  IVSVTX0H U1019 ( .A(n886), .Z(n887) );
  AO7SVTX1 U1020 ( .A(n893), .B(n892), .C(n891), .Z(n895) );
  IVSVTX0H U1021 ( .A(n902), .Z(n903) );
endmodule

