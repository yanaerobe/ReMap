
module m_rangemapping ( N, O );
  input [31:0] N;
  output [31:0] O;
  wire   n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648;

  ND3SVTX1 U296 ( .A(n228), .B(N[1]), .C(n377), .Z(n216) );
  NR3SVTX1 U297 ( .A(n511), .B(n534), .C(n542), .Z(n510) );
  ND3SVTX1 U298 ( .A(N[21]), .B(n226), .C(n268), .Z(n222) );
  ND2SVTX1 U299 ( .A(n235), .B(n263), .Z(n215) );
  ND2SVTX1 U300 ( .A(n236), .B(n244), .Z(n217) );
  NR4SVTX1 U301 ( .A(N[15]), .B(N[14]), .C(N[12]), .D(N[13]), .Z(n236) );
  AO20SVTX1 U302 ( .A(n534), .B(n542), .C(n511), .D(n510), .Z(n512) );
  NR4SVTX1 U303 ( .A(N[28]), .B(N[31]), .C(N[30]), .D(N[29]), .Z(n235) );
  NR4SVTX1 U304 ( .A(N[24]), .B(N[25]), .C(N[27]), .D(n215), .Z(n226) );
  AO17SVTX1 U305 ( .A(n241), .B(N[19]), .C(N[23]), .D(n226), .Z(n212) );
  NR4SVTX1 U306 ( .A(N[23]), .B(N[22]), .C(N[20]), .D(N[21]), .Z(n241) );
  OR4SVTX1 U307 ( .A(N[7]), .B(N[6]), .C(N[4]), .D(N[5]), .Z(n237) );
  NR4SVTX1 U308 ( .A(N[8]), .B(N[9]), .C(N[10]), .D(N[11]), .Z(n244) );
  NR3SVTX1 U309 ( .A(n243), .B(N[26]), .C(n242), .Z(n249) );
  OR3SVTX1 U310 ( .A(N[25]), .B(N[24]), .C(N[27]), .Z(n242) );
  ND4SVTX1 U311 ( .A(n221), .B(n248), .C(n257), .D(n253), .Z(O[31]) );
  IVSVTX0H U312 ( .A(n217), .Z(n238) );
  NR2ASVTX1 U313 ( .A(n238), .B(n237), .Z(n228) );
  AO2NSVTX1 U314 ( .A(n238), .B(N[7]), .C(n228), .D(N[3]), .Z(n211) );
  AO1SVTX1 U315 ( .A(n236), .B(N[11]), .C(N[15]), .D(n211), .Z(n213) );
  IVSVTX0H U316 ( .A(N[26]), .Z(n263) );
  IVSVTX0H U317 ( .A(n226), .Z(n240) );
  NR2ASVTX1 U318 ( .A(n241), .B(n240), .Z(n230) );
  NR2ASVTX1 U319 ( .A(n230), .B(N[18]), .Z(n221) );
  IVSVTX0H U320 ( .A(N[19]), .Z(n248) );
  IVSVTX0H U321 ( .A(N[16]), .Z(n257) );
  IVSVTX0H U322 ( .A(N[17]), .Z(n253) );
  AO7SVTX1 U323 ( .A(n213), .B(O[31]), .C(n212), .Z(n214) );
  AO1SVTX1 U324 ( .A(n235), .B(N[27]), .C(N[31]), .D(n214), .Z(n234) );
  IVSVTX0H U325 ( .A(N[30]), .Z(n231) );
  AO2ASVTX1 U326 ( .C(N[29]), .D(n231), .A(n215), .B(N[25]), .Z(n224) );
  IVSVTX0H U327 ( .A(O[31]), .Z(n262) );
  IVSVTX0H U328 ( .A(N[10]), .Z(n324) );
  IVSVTX0H U329 ( .A(N[5]), .Z(n245) );
  IVSVTX0H U330 ( .A(N[2]), .Z(n377) );
  AO21SVTX1 U331 ( .A(N[6]), .B(n217), .C(n245), .D(n216), .Z(n218) );
  AO8SVTX1 U332 ( .A(n236), .B(N[9]), .C(n324), .D(n218), .Z(n219) );
  AO7ASVTX1 U333 ( .A(N[13]), .B(N[14]), .C(n219), .Z(n220) );
  AO2SVTX1 U334 ( .A(N[17]), .B(n221), .C(n262), .D(n220), .Z(n223) );
  IVSVTX0H U335 ( .A(N[22]), .Z(n268) );
  ND4SVTX1 U336 ( .A(n234), .B(n224), .C(n223), .D(n222), .Z(n225) );
  IVSVTX1 U337 ( .A(n225), .Z(n397) );
  IVSVTX1 U338 ( .A(n397), .Z(O[27]) );
  AO2SVTX1 U339 ( .A(N[22]), .B(n226), .C(N[26]), .D(n235), .Z(n233) );
  AO17NSVTX1 U340 ( .A(n244), .B(N[6]), .C(N[10]), .D(n236), .Z(n227) );
  AO1NSVTX1 U341 ( .A(n228), .B(N[2]), .C(n227), .D(N[14]), .Z(n229) );
  AO2SVTX1 U342 ( .A(n230), .B(N[18]), .C(n262), .D(n229), .Z(n232) );
  ND4SVTX1 U343 ( .A(n234), .B(n233), .C(n232), .D(n231), .Z(O[28]) );
  AO7SVTX1 U344 ( .A(n236), .B(O[31]), .C(n235), .Z(n243) );
  AO8SVTX1 U345 ( .A(n262), .B(n238), .C(n237), .D(n243), .Z(n239) );
  AO7SVTX1 U346 ( .A(n241), .B(n240), .C(n239), .Z(O[29]) );
  AO7SVTX1 U347 ( .A(n244), .B(O[31]), .C(n249), .Z(O[30]) );
  NR2ASVTX1 U348 ( .A(O[30]), .B(O[31]), .Z(n297) );
  AO20CSVTX1 U349 ( .A(O[31]), .B(n245), .C(N[21]), .D(O[30]), .Z(n246) );
  AO1SVTX1 U350 ( .A(N[13]), .B(n297), .C(N[29]), .D(n246), .Z(n256) );
  IVSVTX1 U351 ( .A(O[28]), .Z(n373) );
  NR2ASVTX1 U352 ( .A(O[29]), .B(n373), .Z(n354) );
  IVSVTX0H U353 ( .A(n354), .Z(n339) );
  NR2SVTX1 U354 ( .A(n262), .B(n249), .Z(n363) );
  NR2ASVTX1 U355 ( .A(n363), .B(O[29]), .Z(n367) );
  IVSVTX0H U356 ( .A(O[29]), .Z(n362) );
  IVSVTX0H U357 ( .A(O[30]), .Z(n261) );
  NR2ASVTX1 U358 ( .A(n261), .B(O[31]), .Z(n266) );
  AO2SVTX1 U359 ( .A(n262), .B(N[11]), .C(N[3]), .D(n266), .Z(n247) );
  AO7SVTX1 U360 ( .A(n248), .B(O[30]), .C(n247), .Z(n251) );
  NR2ASVTX1 U361 ( .A(n249), .B(n262), .Z(n342) );
  AO2SVTX1 U362 ( .A(N[15]), .B(n342), .C(N[7]), .D(n297), .Z(n292) );
  IVSVTX0H U363 ( .A(n292), .Z(n250) );
  AO35SVTX1 U364 ( .A(n362), .B(N[27]), .C(n251), .D(O[29]), .E(n250), .Z(n252) );
  AO7ABSVTX1 U365 ( .A(N[23]), .B(n367), .C(n252), .Z(n275) );
  IVSVTX0H U366 ( .A(N[1]), .Z(n468) );
  AO20SVTX1 U367 ( .A(O[31]), .B(n468), .C(n253), .D(O[30]), .Z(n254) );
  AO1SVTX1 U368 ( .A(n262), .B(N[9]), .C(N[25]), .D(n254), .Z(n286) );
  NR2ASVTX1 U369 ( .A(n362), .B(n373), .Z(n348) );
  AO2ASVTX1 U370 ( .C(n373), .D(n275), .A(n286), .B(n348), .Z(n255) );
  AO7SVTX1 U371 ( .A(n256), .B(n339), .C(n255), .Z(n274) );
  BFSVTX1 U372 ( .A(n397), .Z(n470) );
  IVSVTX0H U373 ( .A(N[0]), .Z(n469) );
  AO20SVTX1 U374 ( .A(O[31]), .B(n469), .C(n257), .D(O[30]), .Z(n258) );
  AO1SVTX1 U375 ( .A(n262), .B(N[8]), .C(N[24]), .D(n258), .Z(n278) );
  AO2SVTX1 U376 ( .A(N[20]), .B(n342), .C(N[4]), .D(n266), .Z(n259) );
  AO7SVTX1 U377 ( .A(n278), .B(O[29]), .C(n259), .Z(n260) );
  AO1SVTX1 U378 ( .A(N[12]), .B(n297), .C(N[28]), .D(n260), .Z(n272) );
  AO17SVTX1 U379 ( .A(n262), .B(N[2]), .C(N[18]), .D(n261), .Z(n264) );
  AO3SVTX1 U380 ( .A(O[31]), .B(n324), .C(n264), .D(n263), .Z(n279) );
  NR2ASVTX1 U381 ( .A(O[29]), .B(O[28]), .Z(n337) );
  AO4ABSVTX1 U382 ( .C(n373), .D(n272), .A(n279), .B(n337), .Z(n277) );
  NR2ASVTX1 U383 ( .A(n362), .B(O[28]), .Z(n328) );
  ND2SVTX1 U384 ( .A(n328), .B(n470), .Z(n390) );
  AO11SVTX1 U385 ( .A(N[22]), .B(n363), .C(N[6]), .D(n297), .E(n342), .F(N[14]), .Z(n281) );
  IVSVTX0H U386 ( .A(n281), .Z(n295) );
  AO2ASVTX1 U387 ( .C(n470), .D(n277), .A(n390), .B(n295), .Z(n265) );
  AO7ASVTX1 U388 ( .A(n274), .B(n470), .C(n265), .Z(n498) );
  AO2SVTX1 U389 ( .A(N[14]), .B(n297), .C(N[6]), .D(n266), .Z(n271) );
  IVSVTX0H U390 ( .A(n342), .Z(n322) );
  AO7SVTX1 U392 ( .A(n268), .B(n322), .C(1'b1), .Z(n269) );
  AO1SVTX1 U393 ( .A(n348), .B(n279), .C(N[30]), .D(n269), .Z(n270) );
  AO3SVTX1 U394 ( .A(n272), .B(O[28]), .C(n271), .D(n270), .Z(n273) );
  AO7SVTX1 U395 ( .A(n274), .B(O[27]), .C(n273), .Z(n528) );
  NR2ASVTX1 U396 ( .A(n498), .B(n528), .Z(n642) );
  IVSVTX0H U397 ( .A(n337), .Z(n325) );
  AO4ABSVTX1 U398 ( .C(n286), .D(n325), .A(O[28]), .B(n275), .Z(n283) );
  ND2SVTX1 U399 ( .A(n328), .B(O[27]), .Z(n392) );
  AO11SVTX1 U400 ( .A(N[21]), .B(n363), .C(N[13]), .D(n342), .E(N[5]), .F(n297), .Z(n300) );
  AO4SVTX1 U401 ( .A(n281), .B(n392), .C(n300), .D(n390), .Z(n276) );
  AO10SVTX1 U402 ( .A(n397), .B(n283), .C(O[27]), .D(n277), .E(n276), .Z(n491)
         );
  IVSVTX1 U403 ( .A(n348), .Z(n356) );
  IVSVTX0H U404 ( .A(n278), .Z(n284) );
  AO2SVTX1 U405 ( .A(n354), .B(n279), .C(n337), .D(n284), .Z(n280) );
  AO7SVTX1 U406 ( .A(n281), .B(n356), .C(n280), .Z(n395) );
  AO11SVTX1 U407 ( .A(N[20]), .B(n363), .C(N[12]), .D(n342), .E(N[4]), .F(n297), .Z(n393) );
  AO4SVTX1 U408 ( .A(n300), .B(n392), .C(n393), .D(n390), .Z(n282) );
  AO10SVTX1 U409 ( .A(n397), .B(n395), .C(n225), .D(n283), .E(n282), .Z(n499)
         );
  IVSVTX0H U410 ( .A(n499), .Z(n487) );
  AO2SVTX1 U411 ( .A(n354), .B(n284), .C(n337), .D(n295), .Z(n285) );
  AO7SVTX1 U412 ( .A(n393), .B(n356), .C(n285), .Z(n294) );
  IVSVTX0H U413 ( .A(n363), .Z(n323) );
  NR2ASVTX1 U414 ( .A(n337), .B(n323), .Z(n370) );
  AO4SVTX1 U415 ( .A(n286), .B(n339), .C(n300), .D(n356), .Z(n287) );
  AO6SVTX1 U416 ( .A(N[23]), .B(n370), .C(n287), .Z(n288) );
  AO7SVTX1 U417 ( .A(n292), .B(n325), .C(n288), .Z(n396) );
  AO11SVTX1 U418 ( .A(N[18]), .B(n363), .C(N[10]), .D(n342), .E(N[2]), .F(n297), .Z(n304) );
  AO11SVTX1 U419 ( .A(N[19]), .B(n363), .C(N[11]), .D(n342), .E(N[3]), .F(n297), .Z(n391) );
  AO4SVTX1 U420 ( .A(n304), .B(n390), .C(n391), .D(n392), .Z(n289) );
  AO10SVTX1 U421 ( .A(n397), .B(n294), .C(O[27]), .D(n396), .E(n289), .Z(n495)
         );
  NR2SVTX1 U422 ( .A(n323), .B(n339), .Z(n471) );
  AO4SVTX1 U423 ( .A(n300), .B(n325), .C(n391), .D(n356), .Z(n290) );
  AO6SVTX1 U424 ( .A(N[23]), .B(n471), .C(n290), .Z(n291) );
  AO7SVTX1 U425 ( .A(n292), .B(n339), .C(n291), .Z(n299) );
  AO11SVTX1 U426 ( .A(N[17]), .B(n363), .C(N[9]), .D(n342), .E(N[1]), .F(n297), 
        .Z(n317) );
  AO4SVTX1 U427 ( .A(n304), .B(n392), .C(n317), .D(n390), .Z(n293) );
  AO10SVTX1 U428 ( .A(n397), .B(n299), .C(O[27]), .D(n294), .E(n293), .Z(n515)
         );
  IVSVTX0H U429 ( .A(n393), .Z(n305) );
  AO2SVTX1 U430 ( .A(n354), .B(n295), .C(n337), .D(n305), .Z(n296) );
  AO7SVTX1 U431 ( .A(n304), .B(n356), .C(n296), .Z(n303) );
  AO11SVTX1 U432 ( .A(N[16]), .B(n363), .C(N[8]), .D(n342), .E(n297), .F(N[0]), 
        .Z(n326) );
  AO4SVTX1 U433 ( .A(n317), .B(n392), .C(n326), .D(n390), .Z(n298) );
  AO10SVTX1 U434 ( .A(n397), .B(n303), .C(O[27]), .D(n299), .E(n298), .Z(n520)
         );
  IVSVTX0H U435 ( .A(n391), .Z(n309) );
  AO2ASVTX1 U436 ( .C(n337), .D(n309), .A(n300), .B(n354), .Z(n301) );
  AO7SVTX1 U437 ( .A(n317), .B(n356), .C(n301), .Z(n308) );
  AO2SVTX1 U438 ( .A(N[15]), .B(n363), .C(N[7]), .D(n342), .Z(n331) );
  AO4SVTX1 U439 ( .A(n326), .B(n392), .C(n331), .D(n390), .Z(n302) );
  AO10SVTX1 U440 ( .A(n397), .B(n308), .C(n225), .D(n303), .E(n302), .Z(n526)
         );
  IVSVTX0H U441 ( .A(n304), .Z(n313) );
  AO2SVTX1 U442 ( .A(n354), .B(n305), .C(n337), .D(n313), .Z(n306) );
  AO7SVTX1 U443 ( .A(n326), .B(n356), .C(n306), .Z(n312) );
  AO2SVTX1 U444 ( .A(N[14]), .B(n363), .C(N[6]), .D(n342), .Z(n340) );
  AO4SVTX1 U445 ( .A(n331), .B(n392), .C(n340), .D(n390), .Z(n307) );
  AO10SVTX1 U446 ( .A(n470), .B(n312), .C(O[27]), .D(n308), .E(n307), .Z(n530)
         );
  AO2ASVTX1 U447 ( .C(n354), .D(n309), .A(n317), .B(n337), .Z(n310) );
  AO7SVTX1 U448 ( .A(n331), .B(n356), .C(n310), .Z(n316) );
  AO2SVTX1 U449 ( .A(N[13]), .B(n363), .C(N[5]), .D(n342), .Z(n332) );
  AO4SVTX1 U450 ( .A(n340), .B(n392), .C(n332), .D(n390), .Z(n311) );
  AO10SVTX1 U451 ( .A(n470), .B(n316), .C(n225), .D(n312), .E(n311), .Z(n570)
         );
  AO2ASVTX1 U452 ( .C(n354), .D(n313), .A(n326), .B(n337), .Z(n314) );
  AO7SVTX1 U453 ( .A(n340), .B(n356), .C(n314), .Z(n321) );
  AO2SVTX1 U454 ( .A(N[12]), .B(n363), .C(N[4]), .D(n342), .Z(n336) );
  AO4SVTX1 U455 ( .A(n332), .B(n392), .C(n336), .D(n390), .Z(n315) );
  AO10SVTX1 U456 ( .A(n470), .B(n321), .C(n225), .D(n316), .E(n315), .Z(n574)
         );
  AO2NSVTX1 U457 ( .A(N[11]), .B(n363), .C(N[3]), .D(n342), .Z(n345) );
  AO4SVTX1 U458 ( .A(n317), .B(n339), .C(n331), .D(n325), .Z(n318) );
  AO6SVTX1 U459 ( .A(n328), .B(n345), .C(n318), .Z(n319) );
  AO7SVTX1 U460 ( .A(n332), .B(n356), .C(n319), .Z(n330) );
  NR2SVTX1 U461 ( .A(n336), .B(n392), .Z(n320) );
  AO10SVTX1 U462 ( .A(n397), .B(n330), .C(n225), .D(n321), .E(n320), .Z(n578)
         );
  AO4SVTX1 U463 ( .A(n324), .B(n323), .C(n377), .D(n322), .Z(n352) );
  AO4SVTX1 U464 ( .A(n326), .B(n339), .C(n340), .D(n325), .Z(n327) );
  AO6SVTX1 U465 ( .A(n328), .B(n352), .C(n327), .Z(n329) );
  AO7SVTX1 U466 ( .A(n336), .B(n356), .C(n329), .Z(n335) );
  AO2SVTX1 U467 ( .A(n470), .B(n335), .C(n330), .D(O[27]), .Z(n582) );
  IVSVTX0H U468 ( .A(n331), .Z(n333) );
  IVSVTX0H U469 ( .A(n332), .Z(n347) );
  AO11SVTX1 U470 ( .A(n345), .B(n348), .C(n333), .D(n354), .E(n347), .F(n337), 
        .Z(n341) );
  AO2SVTX1 U471 ( .A(N[9]), .B(n363), .C(N[1]), .D(n342), .Z(n346) );
  AO4SVTX1 U472 ( .A(n341), .B(n225), .C(n346), .D(n390), .Z(n334) );
  AO6SVTX1 U473 ( .A(n225), .B(n335), .C(n334), .Z(n586) );
  IVSVTX0H U474 ( .A(n336), .Z(n353) );
  AO2SVTX1 U475 ( .A(n348), .B(n352), .C(n337), .D(n353), .Z(n338) );
  AO7SVTX1 U476 ( .A(n340), .B(n339), .C(n338), .Z(n351) );
  IVSVTX0H U477 ( .A(n341), .Z(n344) );
  AO2SVTX1 U478 ( .A(N[8]), .B(n363), .C(n342), .D(N[0]), .Z(n358) );
  AO4SVTX1 U479 ( .A(n346), .B(n392), .C(n358), .D(n390), .Z(n343) );
  AO10SVTX1 U480 ( .A(n470), .B(n351), .C(n225), .D(n344), .E(n343), .Z(n590)
         );
  AO2SVTX1 U481 ( .A(O[29]), .B(n345), .C(N[7]), .D(n367), .Z(n361) );
  IVSVTX0H U482 ( .A(n361), .Z(n349) );
  IVSVTX0H U483 ( .A(n346), .Z(n360) );
  AO11SVTX1 U484 ( .A(n349), .B(n373), .C(n360), .D(n348), .E(n347), .F(n354), 
        .Z(n357) );
  AO4SVTX1 U485 ( .A(n358), .B(n392), .C(n357), .D(n225), .Z(n350) );
  AO6SVTX1 U486 ( .A(n225), .B(n351), .C(n350), .Z(n594) );
  AO2SVTX1 U487 ( .A(O[29]), .B(n352), .C(N[6]), .D(n367), .Z(n359) );
  AO2ASVTX1 U488 ( .C(n354), .D(n353), .A(n359), .B(n373), .Z(n355) );
  AO7SVTX1 U489 ( .A(n358), .B(n356), .C(n355), .Z(n388) );
  AO2ASVTX1 U490 ( .C(n470), .D(n388), .A(n357), .B(n225), .Z(n598) );
  AO2ASVTX1 U491 ( .C(N[4]), .D(n367), .A(n358), .B(O[29]), .Z(n364) );
  AO2SVTX1 U492 ( .A(n373), .B(n364), .C(n359), .D(O[28]), .Z(n386) );
  AO2SVTX1 U493 ( .A(N[5]), .B(n367), .C(O[29]), .D(n360), .Z(n365) );
  AO2SVTX1 U494 ( .A(n373), .B(n365), .C(n361), .D(O[28]), .Z(n389) );
  AO2SVTX1 U495 ( .A(n470), .B(n386), .C(n389), .D(n225), .Z(n606) );
  NR2ASVTX1 U496 ( .A(n363), .B(n362), .Z(n368) );
  AO2SVTX1 U497 ( .A(N[6]), .B(n368), .C(N[2]), .D(n367), .Z(n366) );
  AO2SVTX1 U498 ( .A(n373), .B(n366), .C(n364), .D(O[28]), .Z(n384) );
  AO2SVTX1 U499 ( .A(N[7]), .B(n368), .C(N[3]), .D(n367), .Z(n369) );
  AO2SVTX1 U500 ( .A(n373), .B(n369), .C(n365), .D(O[28]), .Z(n387) );
  AO2SVTX1 U501 ( .A(n470), .B(n384), .C(n387), .D(n225), .Z(n614) );
  AO2SVTX1 U502 ( .A(N[4]), .B(n368), .C(n367), .D(N[0]), .Z(n371) );
  AO2SVTX1 U503 ( .A(n373), .B(n371), .C(n366), .D(O[28]), .Z(n382) );
  AO2SVTX1 U504 ( .A(N[5]), .B(n368), .C(N[1]), .D(n367), .Z(n372) );
  AO2SVTX1 U505 ( .A(n373), .B(n372), .C(n369), .D(O[28]), .Z(n385) );
  AO2SVTX1 U506 ( .A(n470), .B(n382), .C(n385), .D(O[27]), .Z(n622) );
  IVSVTX0H U507 ( .A(n370), .Z(n376) );
  AO4SVTX1 U508 ( .A(n373), .B(n371), .C(n377), .D(n376), .Z(n375) );
  IVSVTX0H U509 ( .A(N[3]), .Z(n374) );
  AO4SVTX1 U510 ( .A(n373), .B(n372), .C(n374), .D(n376), .Z(n383) );
  AO2SVTX1 U511 ( .A(n470), .B(n375), .C(n383), .D(O[27]), .Z(n630) );
  AO7SVTX1 U512 ( .A(N[1]), .B(N[0]), .C(n471), .Z(n380) );
  IVSVTX0H U513 ( .A(n471), .Z(n467) );
  AO4SVTX1 U514 ( .A(n374), .B(n467), .C(n468), .D(n376), .Z(n378) );
  AO2SVTX1 U515 ( .A(n470), .B(n378), .C(n375), .D(O[27]), .Z(n634) );
  AO4SVTX1 U516 ( .A(n377), .B(n467), .C(n469), .D(n376), .Z(n379) );
  AO2SVTX1 U517 ( .A(n470), .B(n379), .C(n378), .D(O[27]), .Z(n484) );
  AO9SVTX1 U518 ( .A(N[1]), .B(n397), .C(n471), .D(n379), .E(O[27]), .Z(n474)
         );
  ND4SVTX1 U519 ( .A(n380), .B(n634), .C(n484), .D(n474), .Z(n381) );
  NR2ASVTX1 U520 ( .A(n630), .B(n381), .Z(n462) );
  AO2SVTX1 U521 ( .A(n470), .B(n383), .C(n382), .D(O[27]), .Z(n626) );
  ND2SVTX1 U522 ( .A(n462), .B(n626), .Z(n461) );
  NR2ASVTX1 U523 ( .A(n622), .B(n461), .Z(n458) );
  AO2SVTX1 U524 ( .A(n470), .B(n385), .C(n384), .D(O[27]), .Z(n618) );
  ND2SVTX1 U525 ( .A(n458), .B(n618), .Z(n455) );
  NR2ASVTX1 U526 ( .A(n614), .B(n455), .Z(n452) );
  AO2SVTX1 U527 ( .A(n470), .B(n387), .C(n386), .D(O[27]), .Z(n610) );
  ND2SVTX1 U528 ( .A(n452), .B(n610), .Z(n449) );
  NR2ASVTX1 U529 ( .A(n606), .B(n449), .Z(n446) );
  AO2SVTX1 U530 ( .A(n470), .B(n389), .C(n388), .D(O[27]), .Z(n602) );
  ND2SVTX1 U531 ( .A(n446), .B(n602), .Z(n443) );
  NR2ASVTX1 U532 ( .A(n598), .B(n443), .Z(n440) );
  ND2SVTX1 U533 ( .A(n594), .B(n440), .Z(n437) );
  NR2ASVTX1 U534 ( .A(n590), .B(n437), .Z(n434) );
  ND2SVTX1 U535 ( .A(n586), .B(n434), .Z(n431) );
  NR2ASVTX1 U536 ( .A(n582), .B(n431), .Z(n428) );
  ND2SVTX1 U537 ( .A(n578), .B(n428), .Z(n425) );
  NR2ASVTX1 U538 ( .A(n574), .B(n425), .Z(n422) );
  ND2SVTX1 U539 ( .A(n570), .B(n422), .Z(n419) );
  NR2ASVTX1 U540 ( .A(n530), .B(n419), .Z(n416) );
  ND2SVTX1 U541 ( .A(n526), .B(n416), .Z(n413) );
  NR2ASVTX1 U542 ( .A(n520), .B(n413), .Z(n410) );
  ND2SVTX1 U543 ( .A(n515), .B(n410), .Z(n407) );
  NR2ASVTX1 U544 ( .A(n495), .B(n407), .Z(n404) );
  AO4SVTX1 U545 ( .A(n393), .B(n392), .C(n391), .D(n390), .Z(n394) );
  AO10SVTX1 U546 ( .A(n397), .B(n396), .C(O[27]), .D(n395), .E(n394), .Z(n489)
         );
  ND2SVTX1 U547 ( .A(n404), .B(n489), .Z(n401) );
  NR2ASVTX1 U548 ( .A(n499), .B(n401), .Z(n399) );
  ND2SVTX1 U549 ( .A(n491), .B(n399), .Z(n500) );
  NR2SVTX1 U550 ( .A(n528), .B(n498), .Z(n504) );
  BFSVTX1 U551 ( .A(n642), .Z(n479) );
  AO7NSVTX1 U552 ( .A(n491), .B(n399), .C(n500), .Z(n400) );
  IVSVTX0H U553 ( .A(n491), .Z(n398) );
  NR2ASVTX1 U554 ( .A(n528), .B(n498), .Z(n641) );
  IVSVTX0H U555 ( .A(n641), .Z(n645) );
  IVSVTX1 U556 ( .A(n645), .Z(n507) );
  AO11SVTX1 U557 ( .A(n500), .B(n504), .C(n479), .D(n400), .E(n398), .F(n507), 
        .Z(n490) );
  AO6SVTX1 U558 ( .A(n487), .B(n401), .C(n399), .Z(n402) );
  AO11SVTX1 U559 ( .A(n487), .B(n507), .C(n479), .D(n402), .E(n400), .F(n504), 
        .Z(n496) );
  IVSVTX0H U560 ( .A(n489), .Z(n403) );
  AO7NSVTX1 U561 ( .A(n404), .B(n489), .C(n401), .Z(n405) );
  AO11SVTX1 U562 ( .A(n403), .B(n641), .C(n504), .D(n402), .E(n479), .F(n405), 
        .Z(n516) );
  IVSVTX0H U563 ( .A(n495), .Z(n406) );
  AO6SVTX1 U564 ( .A(n406), .B(n407), .C(n404), .Z(n408) );
  AO11SVTX1 U565 ( .A(n406), .B(n641), .C(n504), .D(n405), .E(n642), .F(n408), 
        .Z(n521) );
  IVSVTX0H U566 ( .A(n515), .Z(n409) );
  AO7NSVTX1 U567 ( .A(n515), .B(n410), .C(n407), .Z(n411) );
  AO11SVTX1 U568 ( .A(n409), .B(n641), .C(n504), .D(n408), .E(n642), .F(n411), 
        .Z(n527) );
  IVSVTX0H U569 ( .A(n520), .Z(n412) );
  AO6SVTX1 U570 ( .A(n412), .B(n413), .C(n410), .Z(n414) );
  AO11SVTX1 U571 ( .A(n412), .B(n641), .C(n504), .D(n411), .E(n642), .F(n414), 
        .Z(n531) );
  IVSVTX0H U572 ( .A(n526), .Z(n415) );
  AO7NSVTX1 U573 ( .A(n526), .B(n416), .C(n413), .Z(n417) );
  AO11SVTX1 U574 ( .A(n415), .B(n507), .C(n504), .D(n414), .E(n479), .F(n417), 
        .Z(n571) );
  IVSVTX0H U575 ( .A(n530), .Z(n418) );
  AO6SVTX1 U576 ( .A(n418), .B(n419), .C(n416), .Z(n420) );
  AO11SVTX1 U577 ( .A(n418), .B(n507), .C(n504), .D(n417), .E(n642), .F(n420), 
        .Z(n575) );
  IVSVTX0H U578 ( .A(n570), .Z(n421) );
  BFSVTX1 U579 ( .A(n504), .Z(n493) );
  AO7NSVTX1 U580 ( .A(n570), .B(n422), .C(n419), .Z(n423) );
  AO11SVTX1 U581 ( .A(n421), .B(n507), .C(n493), .D(n420), .E(n479), .F(n423), 
        .Z(n579) );
  IVSVTX0H U582 ( .A(n574), .Z(n424) );
  AO6SVTX1 U583 ( .A(n424), .B(n425), .C(n422), .Z(n426) );
  AO11SVTX1 U584 ( .A(n424), .B(n507), .C(n493), .D(n423), .E(n642), .F(n426), 
        .Z(n583) );
  IVSVTX0H U585 ( .A(n578), .Z(n427) );
  AO7NSVTX1 U586 ( .A(n578), .B(n428), .C(n425), .Z(n430) );
  AO11SVTX1 U587 ( .A(n427), .B(n507), .C(n493), .D(n426), .E(n479), .F(n430), 
        .Z(n587) );
  IVSVTX0H U588 ( .A(n582), .Z(n429) );
  AO6SVTX1 U589 ( .A(n429), .B(n431), .C(n428), .Z(n432) );
  AO11SVTX1 U590 ( .A(n642), .B(n432), .C(n493), .D(n430), .E(n429), .F(n507), 
        .Z(n591) );
  IVSVTX0H U591 ( .A(n586), .Z(n433) );
  AO7NSVTX1 U592 ( .A(n586), .B(n434), .C(n431), .Z(n435) );
  AO11SVTX1 U593 ( .A(n433), .B(n507), .C(n493), .D(n432), .E(n479), .F(n435), 
        .Z(n595) );
  IVSVTX0H U594 ( .A(n590), .Z(n436) );
  AO6SVTX1 U595 ( .A(n436), .B(n437), .C(n434), .Z(n438) );
  AO11SVTX1 U596 ( .A(n436), .B(n507), .C(n493), .D(n435), .E(n479), .F(n438), 
        .Z(n599) );
  IVSVTX0H U597 ( .A(n594), .Z(n439) );
  AO7NSVTX1 U598 ( .A(n594), .B(n440), .C(n437), .Z(n442) );
  AO11SVTX1 U599 ( .A(n439), .B(n507), .C(n493), .D(n438), .E(n479), .F(n442), 
        .Z(n603) );
  IVSVTX0H U600 ( .A(n598), .Z(n441) );
  AO6SVTX1 U601 ( .A(n441), .B(n443), .C(n440), .Z(n445) );
  AO11SVTX1 U602 ( .A(n642), .B(n445), .C(n493), .D(n442), .E(n441), .F(n507), 
        .Z(n607) );
  AO7NSVTX1 U603 ( .A(n446), .B(n602), .C(n443), .Z(n448) );
  IVSVTX0H U604 ( .A(n602), .Z(n444) );
  AO11SVTX1 U605 ( .A(n479), .B(n448), .C(n493), .D(n445), .E(n444), .F(n507), 
        .Z(n611) );
  IVSVTX0H U606 ( .A(n606), .Z(n447) );
  AO6SVTX1 U607 ( .A(n447), .B(n449), .C(n446), .Z(n451) );
  AO11SVTX1 U608 ( .A(n479), .B(n451), .C(n493), .D(n448), .E(n447), .F(n507), 
        .Z(n615) );
  AO7NSVTX1 U609 ( .A(n452), .B(n610), .C(n449), .Z(n454) );
  IVSVTX0H U610 ( .A(n610), .Z(n450) );
  AO11SVTX1 U611 ( .A(n479), .B(n454), .C(n493), .D(n451), .E(n450), .F(n507), 
        .Z(n619) );
  IVSVTX0H U612 ( .A(n614), .Z(n453) );
  AO6SVTX1 U613 ( .A(n453), .B(n455), .C(n452), .Z(n457) );
  AO11SVTX1 U614 ( .A(n479), .B(n457), .C(n493), .D(n454), .E(n453), .F(n507), 
        .Z(n623) );
  AO7NSVTX1 U615 ( .A(n458), .B(n618), .C(n455), .Z(n460) );
  IVSVTX0H U616 ( .A(n618), .Z(n456) );
  AO11SVTX1 U617 ( .A(n479), .B(n460), .C(n493), .D(n457), .E(n456), .F(n507), 
        .Z(n627) );
  IVSVTX0H U618 ( .A(n622), .Z(n459) );
  AO6SVTX1 U619 ( .A(n459), .B(n461), .C(n458), .Z(n464) );
  AO11SVTX1 U620 ( .A(n479), .B(n464), .C(n493), .D(n460), .E(n459), .F(n507), 
        .Z(n631) );
  AO7NSVTX1 U621 ( .A(n462), .B(n626), .C(n461), .Z(n465) );
  IVSVTX0H U622 ( .A(n626), .Z(n463) );
  AO11SVTX1 U623 ( .A(n479), .B(n465), .C(n493), .D(n464), .E(n463), .F(n507), 
        .Z(n635) );
  AO4ABSVTX1 U624 ( .C(n630), .D(n645), .A(n493), .B(n465), .Z(n466) );
  AO6SVTX1 U625 ( .A(n479), .B(n630), .C(n466), .Z(n486) );
  IVSVTX0H U626 ( .A(n474), .Z(n483) );
  AO10SVTX1 U627 ( .A(n470), .B(n469), .C(O[27]), .D(n468), .E(n467), .Z(n478)
         );
  AO2SVTX1 U628 ( .A(n479), .B(n474), .C(n493), .D(n484), .Z(n473) );
  ND3SVTX1 U629 ( .A(N[0]), .B(n471), .C(O[27]), .Z(n472) );
  AO20SVTX1 U630 ( .A(n474), .B(n645), .C(n473), .D(n472), .Z(n477) );
  AO2SVTX1 U631 ( .A(n479), .B(n484), .C(n493), .D(n634), .Z(n475) );
  AO7SVTX1 U632 ( .A(n484), .B(n645), .C(n475), .Z(n476) );
  AO5NSVTX1 U633 ( .A(n478), .B(n477), .C(n476), .Z(n482) );
  AO2SVTX1 U634 ( .A(n479), .B(n634), .C(n493), .D(n630), .Z(n480) );
  AO7SVTX1 U635 ( .A(n634), .B(n645), .C(n480), .Z(n481) );
  AO5SVTX1 U636 ( .A(n483), .B(n482), .C(n481), .Z(n485) );
  FA1SVTX1 U637 ( .A(n486), .B(n485), .CI(n484), .CO(n633) );
  NR2ASVTX1 U638 ( .A(n487), .B(n502), .Z(n492) );
  NR2ASVTX1 U639 ( .A(n491), .B(n492), .Z(n532) );
  IVSVTX0H U640 ( .A(n532), .Z(n534) );
  FA1SVTX1 U641 ( .A(n490), .B(n489), .CI(n488), .CO(n502), .Z(n546) );
  ND2ASVTX1 U642 ( .A(n546), .B(n532), .Z(n518) );
  NR2ASVTX1 U643 ( .A(n492), .B(n491), .Z(n640) );
  IVSVTX0H U644 ( .A(n640), .Z(n646) );
  AO2SVTX1 U645 ( .A(n493), .B(n646), .C(n528), .D(n534), .Z(n517) );
  FA1SVTX1 U646 ( .A(n496), .B(n495), .CI(n494), .CO(n488), .Z(n550) );
  NR2ASVTX1 U647 ( .A(n646), .B(n532), .Z(n643) );
  ND2SVTX1 U648 ( .A(n498), .B(n528), .Z(n497) );
  AO7SVTX1 U649 ( .A(n643), .B(n528), .C(n497), .Z(n523) );
  ND3ABSVTX1 U650 ( .A(n550), .B(n534), .C(n523), .Z(n522) );
  IVSVTX0H U651 ( .A(n497), .Z(n505) );
  IVSVTX0H U652 ( .A(n643), .Z(n539) );
  AO7SVTX1 U653 ( .A(n498), .B(n539), .C(n646), .Z(n535) );
  AO1SVTX1 U654 ( .A(n532), .B(n505), .C(n504), .D(n535), .Z(n511) );
  AO7SVTX1 U655 ( .A(n528), .B(n500), .C(n499), .Z(n501) );
  EOSVTX1 U656 ( .A(n502), .B(n501), .Z(n542) );
  NR2ASVTX1 U657 ( .A(n513), .B(n510), .Z(n509) );
  AO7SVTX1 U658 ( .A(n642), .B(n534), .C(n509), .Z(n533) );
  MUX21NSVTX1 U659 ( .A(n534), .B(n539), .S(n505), .Z(n503) );
  ND2SVTX1 U660 ( .A(n503), .B(n533), .Z(n637) );
  AO7SVTX1 U661 ( .A(n533), .B(n503), .C(n637), .Z(n543) );
  ND2ASVTX1 U662 ( .A(n533), .B(n532), .Z(n547) );
  NR2ASVTX1 U663 ( .A(n642), .B(n643), .Z(n537) );
  AO20SVTX1 U664 ( .A(n505), .B(n504), .C(n643), .D(n537), .Z(n506) );
  AO7SVTX1 U665 ( .A(n507), .B(n646), .C(n506), .Z(n508) );
  EOSVTX1 U666 ( .A(n509), .B(n508), .Z(n551) );
  EOSVTX1 U667 ( .A(n513), .B(n512), .Z(n555) );
  FA1SVTX1 U668 ( .A(n516), .B(n515), .CI(n514), .CO(n494), .Z(n554) );
  FA1SVTX1 U669 ( .A(n518), .B(n517), .CI(n522), .CO(n513), .Z(n559) );
  FA1SVTX1 U670 ( .A(n521), .B(n520), .CI(n519), .CO(n514), .Z(n558) );
  NR2SVTX1 U671 ( .A(n534), .B(n550), .Z(n524) );
  AO7SVTX1 U672 ( .A(n524), .B(n523), .C(n522), .Z(n563) );
  FA1SVTX1 U673 ( .A(n527), .B(n526), .CI(n525), .CO(n519), .Z(n562) );
  AO2ASVTX1 U674 ( .C(n643), .D(n528), .A(n528), .B(n532), .Z(n567) );
  FA1SVTX1 U675 ( .A(n531), .B(n530), .CI(n529), .CO(n525), .Z(n566) );
  ND2ASVTX1 U676 ( .A(n554), .B(n532), .Z(n565) );
  AO4SVTX1 U677 ( .A(n540), .B(n539), .C(n534), .D(n533), .Z(n638) );
  AO7SVTX1 U678 ( .A(n535), .B(n537), .C(n637), .Z(n536) );
  AO7SVTX1 U679 ( .A(n537), .B(n637), .C(n536), .Z(n639) );
  AO7SVTX1 U680 ( .A(n638), .B(n640), .C(n639), .Z(n538) );
  AO7SVTX1 U681 ( .A(n638), .B(n639), .C(n538), .Z(O[25]) );
  AO6SVTX1 U682 ( .A(n540), .B(n539), .C(n638), .Z(O[24]) );
  FA1SVTX1 U683 ( .A(n543), .B(n542), .CI(n541), .CO(n540), .Z(n544) );
  IVSVTX0H U684 ( .A(n544), .Z(O[23]) );
  FA1SVTX1 U685 ( .A(n547), .B(n546), .CI(n545), .CO(n541), .Z(n548) );
  IVSVTX0H U686 ( .A(n548), .Z(O[22]) );
  FA1SVTX1 U687 ( .A(n551), .B(n550), .CI(n549), .CO(n545), .Z(n552) );
  IVSVTX0H U688 ( .A(n552), .Z(O[21]) );
  FA1SVTX1 U689 ( .A(n555), .B(n554), .CI(n553), .CO(n549), .Z(n556) );
  IVSVTX0H U690 ( .A(n556), .Z(O[20]) );
  FA1SVTX1 U691 ( .A(n559), .B(n558), .CI(n557), .CO(n553), .Z(n560) );
  IVSVTX0H U692 ( .A(n560), .Z(O[19]) );
  FA1SVTX1 U693 ( .A(n563), .B(n562), .CI(n561), .CO(n557), .Z(n564) );
  IVSVTX0H U694 ( .A(n564), .Z(O[18]) );
  FA1SVTX1 U695 ( .A(n567), .B(n566), .CI(n565), .CO(n561), .Z(n568) );
  IVSVTX0H U696 ( .A(n568), .Z(O[17]) );
  FA1SVTX1 U697 ( .A(n571), .B(n570), .CI(n569), .CO(n529), .Z(n572) );
  IVSVTX0H U698 ( .A(n572), .Z(O[16]) );
  FA1SVTX1 U699 ( .A(n575), .B(n574), .CI(n573), .CO(n569), .Z(n576) );
  IVSVTX0H U700 ( .A(n576), .Z(O[15]) );
  FA1SVTX1 U701 ( .A(n579), .B(n578), .CI(n577), .CO(n573), .Z(n580) );
  IVSVTX0H U702 ( .A(n580), .Z(O[14]) );
  FA1SVTX1 U703 ( .A(n583), .B(n582), .CI(n581), .CO(n577), .Z(n584) );
  IVSVTX0H U704 ( .A(n584), .Z(O[13]) );
  FA1SVTX1 U705 ( .A(n587), .B(n586), .CI(n585), .CO(n581), .Z(n588) );
  IVSVTX0H U706 ( .A(n588), .Z(O[12]) );
  FA1SVTX1 U707 ( .A(n591), .B(n590), .CI(n589), .CO(n585), .Z(n592) );
  IVSVTX0H U708 ( .A(n592), .Z(O[11]) );
  FA1SVTX1 U709 ( .A(n595), .B(n594), .CI(n593), .CO(n589), .Z(n596) );
  IVSVTX0H U710 ( .A(n596), .Z(O[10]) );
  FA1SVTX1 U711 ( .A(n599), .B(n598), .CI(n597), .CO(n593), .Z(n600) );
  IVSVTX0H U712 ( .A(n600), .Z(O[9]) );
  FA1SVTX1 U713 ( .A(n603), .B(n602), .CI(n601), .CO(n597), .Z(n604) );
  IVSVTX0H U714 ( .A(n604), .Z(O[8]) );
  FA1SVTX1 U715 ( .A(n607), .B(n606), .CI(n605), .CO(n601), .Z(n608) );
  IVSVTX0H U716 ( .A(n608), .Z(O[7]) );
  FA1SVTX1 U717 ( .A(n611), .B(n610), .CI(n609), .CO(n605), .Z(n612) );
  IVSVTX0H U718 ( .A(n612), .Z(O[6]) );
  FA1SVTX1 U719 ( .A(n615), .B(n614), .CI(n613), .CO(n609), .Z(n616) );
  IVSVTX0H U720 ( .A(n616), .Z(O[5]) );
  FA1SVTX1 U721 ( .A(n619), .B(n618), .CI(n617), .CO(n613), .Z(n620) );
  IVSVTX0H U722 ( .A(n620), .Z(O[4]) );
  FA1SVTX1 U723 ( .A(n623), .B(n622), .CI(n621), .CO(n617), .Z(n624) );
  IVSVTX0H U724 ( .A(n624), .Z(O[3]) );
  FA1SVTX1 U725 ( .A(n627), .B(n626), .CI(n625), .CO(n621), .Z(n628) );
  IVSVTX0H U726 ( .A(n628), .Z(O[2]) );
  FA1SVTX1 U727 ( .A(n631), .B(n630), .CI(n629), .CO(n625), .Z(n632) );
  IVSVTX0H U728 ( .A(n632), .Z(O[1]) );
  FA1SVTX1 U729 ( .A(n635), .B(n634), .CI(n633), .CO(n629), .Z(n636) );
  IVSVTX0H U730 ( .A(n636), .Z(O[0]) );
  AO20DSVTX1 U731 ( .A(n639), .B(n638), .C(n646), .D(n637), .Z(n648) );
  AO1NSVTX1 U732 ( .A(n643), .B(n642), .C(n641), .D(n640), .Z(n644) );
  AO7SVTX1 U733 ( .A(n646), .B(n645), .C(n644), .Z(n647) );
  EOSVTX1 U734 ( .A(n648), .B(n647), .Z(O[26]) );
endmodule

