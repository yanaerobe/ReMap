
module m_rangemapping ( N, O );
  input [31:0] N;
  output [31:0] O;
  wire   n211, n212, n213, n214, n215, n216, n217, n218, n220, n221, n222,
         n223, n225, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n307, n308, n309, n310, n311, n312, n314, n317,
         n318, n319, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n370, n371, n372, n373, n374, n375,
         n377, n378, n379, n380, n381, n383, n384, n385, n386, n387, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830;

  BFSVTX0H U296 ( .A(n386), .Z(O[30]) );
  B_ND2SVTX2 U297 ( .A(n1826), .B(n869), .Z(n1829) );
  IVSVTX0H U298 ( .A(n1721), .Z(n1723) );
  IVSVTX0H U299 ( .A(n1808), .Z(n1810) );
  IVSVTX0H U300 ( .A(n1800), .Z(n1802) );
  IVSVTX0H U301 ( .A(n1713), .Z(n1748) );
  IVSVTX0H U302 ( .A(n1778), .Z(n1779) );
  BFSVTX4 U303 ( .A(n1676), .Z(n810) );
  IVSVTX0H U304 ( .A(n1816), .Z(n1796) );
  IVSVTX0H U305 ( .A(n406), .Z(n1789) );
  IVSVTX0H U306 ( .A(n370), .Z(n1717) );
  IVSVTX0H U307 ( .A(n1787), .Z(n1418) );
  NR2SVTX2 U308 ( .A(n1671), .B(n1670), .Z(n1827) );
  AO7SVTX6 U309 ( .A(n1650), .B(n1649), .C(n1674), .Z(n1651) );
  IVSVTX0H U310 ( .A(n606), .Z(n1792) );
  IVSVTX0H U311 ( .A(n1724), .Z(n1725) );
  IVSVTX0H U312 ( .A(n1781), .Z(n1782) );
  IVSVTX0H U313 ( .A(n1811), .Z(n1812) );
  BFSVTX0H U314 ( .A(n607), .Z(n606) );
  BFSVTX0H U315 ( .A(n1737), .Z(n396) );
  IVSVTX8 U316 ( .A(n525), .Z(n1713) );
  BFSVTX2 U317 ( .A(n1735), .Z(n1742) );
  ND2SVTX6 U318 ( .A(n1646), .B(n1647), .Z(n1680) );
  AO2SVTX2 U319 ( .A(n819), .B(n1665), .C(n1664), .D(n1663), .Z(n1666) );
  AO7ABSVTX6 U320 ( .A(n1635), .B(n1634), .C(n484), .Z(n1639) );
  NR2ASVTX2 U321 ( .A(n1565), .B(n861), .Z(n472) );
  AO7ASVTX6 U322 ( .A(n1626), .B(n1664), .C(n279), .Z(n455) );
  FAS1SVTX2 U323 ( .A(n1580), .B(n280), .CI(n1579), .CO(n1583), .Z(n1633) );
  AN2BSVTX4 U324 ( .A(n1610), .B(n1624), .Z(n1708) );
  ENSVTX0H U325 ( .A(n1550), .B(n1218), .Z(n1242) );
  F_IVSVTX1 U326 ( .A(n1638), .Z(n275) );
  ND2ASVTX6 U327 ( .A(n1601), .B(n861), .Z(n432) );
  NR2SVTX2 U328 ( .A(n1635), .B(n1634), .Z(n486) );
  ND2SVTX2 U329 ( .A(n745), .B(n274), .Z(n478) );
  ND2ASVTX4 U330 ( .A(n1213), .B(n338), .Z(n1560) );
  IVSVTX2 U331 ( .A(n242), .Z(n223) );
  BFSVTX4 U332 ( .A(n474), .Z(n338) );
  IVSVTX0H U333 ( .A(n1578), .Z(n817) );
  BFSVTX4 U334 ( .A(n805), .Z(n802) );
  BFSVTX10 U335 ( .A(n1627), .Z(n1664) );
  BFSVTX0H U336 ( .A(n1605), .Z(n229) );
  IVSVTX2 U337 ( .A(n1581), .Z(n279) );
  IVSVTX0H U338 ( .A(n1616), .Z(n852) );
  IVSVTX6 U339 ( .A(n474), .Z(n274) );
  BFSVTX2 U340 ( .A(n1596), .Z(n241) );
  ND2SVTX2 U341 ( .A(n1620), .B(n1574), .Z(n1576) );
  ND2ASVTX6 U342 ( .A(n395), .B(n1620), .Z(n760) );
  IVSVTX2 U343 ( .A(n1626), .Z(n1601) );
  IVSVTX1 U344 ( .A(n1618), .Z(n1572) );
  IVSVTX0H U345 ( .A(n1212), .Z(n267) );
  NR3SVTX4 U346 ( .A(n748), .B(n1607), .C(n395), .Z(n789) );
  BFSVTX6 U347 ( .A(n1570), .Z(n395) );
  NR2SVTX4 U348 ( .A(n847), .B(n441), .Z(n340) );
  BFSVTX4 U349 ( .A(n1545), .Z(n1619) );
  IVSVTX6 U350 ( .A(n1607), .Z(n1620) );
  ND2ASVTX4 U351 ( .A(n1237), .B(n368), .Z(n1546) );
  CTIVSVTX2 U352 ( .A(n1570), .Z(n713) );
  ND2SVTX6 U353 ( .A(n856), .B(n1618), .Z(n1302) );
  NR2SVTX4 U354 ( .A(n1303), .B(n1305), .Z(n787) );
  ND2ASVTX6 U355 ( .A(n622), .B(n1569), .Z(n1605) );
  ND2ASVTX6 U356 ( .A(n1550), .B(n708), .Z(n856) );
  NR2SVTX6 U357 ( .A(n1535), .B(n1534), .Z(n1721) );
  ND2SVTX4 U358 ( .A(n276), .B(n1596), .Z(n648) );
  ND3ASVTX6 U359 ( .A(n1233), .B(n623), .C(n624), .Z(n1567) );
  IVSVTX0H U360 ( .A(n280), .Z(n622) );
  IVSVTX0H U361 ( .A(n256), .Z(n578) );
  ND3ASVTX6 U362 ( .A(n1523), .B(n641), .C(n640), .Z(n1710) );
  AO7SVTX6 U363 ( .A(n1800), .B(n1804), .C(n1801), .Z(n1813) );
  BFSVTX0H U364 ( .A(n282), .Z(n393) );
  BFSVTX0H U365 ( .A(n1453), .Z(n1455) );
  ND2ASVTX6 U366 ( .A(n288), .B(n333), .Z(n1781) );
  ND2SVTX4 U367 ( .A(n1457), .B(n566), .Z(n565) );
  ND3ASVTX6 U368 ( .A(n1228), .B(n763), .C(n764), .Z(n596) );
  AO7ABSVTX4 U369 ( .A(n1516), .B(n264), .C(n1454), .Z(n562) );
  IVSVTX2 U370 ( .A(n1488), .Z(n278) );
  NR2SVTX2 U371 ( .A(n257), .B(n660), .Z(n664) );
  IVSVTX0H U372 ( .A(n416), .Z(n1002) );
  ND3SVTX4 U373 ( .A(n519), .B(n1417), .C(n518), .Z(n607) );
  ND2SVTX2 U374 ( .A(n636), .B(n877), .Z(n635) );
  ND3SVTX6 U375 ( .A(n245), .B(n669), .C(n1255), .Z(n358) );
  ND2SVTX4 U376 ( .A(n1244), .B(n698), .Z(n697) );
  ND2SVTX6 U377 ( .A(n745), .B(n754), .Z(n634) );
  AO2SVTX4 U378 ( .A(n248), .B(n1379), .C(n1232), .D(n1457), .Z(n1454) );
  OR2BSVTX4 U379 ( .A(n1213), .B(n261), .Z(n1452) );
  AO6SVTX6 U380 ( .A(n747), .B(n255), .C(n746), .Z(n1226) );
  AO7SVTX6 U381 ( .A(n769), .B(n766), .C(n256), .Z(n763) );
  ND3SVTX4 U382 ( .A(n801), .B(n1255), .C(n1215), .Z(n222) );
  AO8ASVTX4 U383 ( .A(n276), .B(n1293), .C(n638), .D(n639), .Z(n637) );
  B_IVSVTX1 U384 ( .A(n385), .Z(n366) );
  IVSVTX4 U385 ( .A(n1275), .Z(n280) );
  ND4ABSVTX6 U386 ( .A(n257), .B(n253), .C(n245), .D(n1255), .Z(n666) );
  IVSVTX2 U387 ( .A(n1492), .Z(n663) );
  ND2ASVTX6 U388 ( .A(n521), .B(n1398), .Z(n644) );
  BFSVTX0H U389 ( .A(n785), .Z(n416) );
  ND2ASVTX6 U390 ( .A(n1228), .B(n1360), .Z(n1411) );
  IVSVTX2 U391 ( .A(n1292), .Z(n638) );
  NR2ASVTX4 U392 ( .A(n1550), .B(n833), .Z(n1233) );
  IVSVTX4 U393 ( .A(n1280), .Z(n256) );
  IVSVTX0H U394 ( .A(n1401), .Z(n284) );
  IVSVTX1 U395 ( .A(n1298), .Z(n239) );
  ND2SVTX4 U396 ( .A(n1516), .B(n1435), .Z(n772) );
  NR2SVTX2 U397 ( .A(n1491), .B(n1823), .Z(n639) );
  IVSVTX4 U398 ( .A(n766), .Z(n765) );
  NR2SVTX2 U399 ( .A(n1416), .B(n1397), .Z(n518) );
  ND2ASVTX4 U400 ( .A(n573), .B(n1443), .Z(n1444) );
  ND2SVTX6 U401 ( .A(n385), .B(n1520), .Z(n481) );
  NR2SVTX6 U402 ( .A(n255), .B(n581), .Z(n627) );
  ND2SVTX6 U403 ( .A(n1516), .B(n1438), .Z(n552) );
  ND2SVTX1 U404 ( .A(n1310), .B(n1232), .Z(n374) );
  IVSVTX0H U405 ( .A(n517), .Z(n237) );
  ND3SVTX4 U406 ( .A(n859), .B(n1604), .C(n660), .Z(n538) );
  AO1CDSVTX4 U407 ( .A(n420), .B(n591), .C(n1516), .D(n1275), .Z(n372) );
  IVSVTX12 U408 ( .A(n1256), .Z(n1255) );
  NR2ASVTX4 U409 ( .A(n1461), .B(n1823), .Z(n1442) );
  IVSVTX8 U410 ( .A(n1557), .Z(n245) );
  IVSVTX0H U411 ( .A(n262), .Z(n517) );
  IVSVTX4 U412 ( .A(n1237), .Z(n255) );
  IVSVTX4 U413 ( .A(n1491), .Z(n276) );
  CTBUFSVTX2 U414 ( .A(n1267), .Z(n217) );
  AO7SVTX4 U415 ( .A(n542), .B(n1491), .C(n1665), .Z(n1292) );
  IVSVTX1 U416 ( .A(n820), .Z(n521) );
  IVSVTX6 U417 ( .A(n483), .Z(n603) );
  ND2SVTX2 U418 ( .A(n548), .B(n1448), .Z(n1456) );
  IVSVTX4 U419 ( .A(n1232), .Z(n771) );
  ND2ASVTX6 U420 ( .A(n1220), .B(n1219), .Z(n1557) );
  ND3ABSVTX6 U421 ( .A(n289), .B(n1490), .C(n1489), .Z(n1535) );
  BFSVTX0H U422 ( .A(n1392), .Z(n1393) );
  BFSVTX0H U423 ( .A(n1091), .Z(n391) );
  IVSVTX2 U424 ( .A(n282), .Z(n722) );
  IVSVTX2 U425 ( .A(n1533), .Z(n277) );
  IVSVTX0H U426 ( .A(n1447), .Z(n1448) );
  IVSVTX0H U427 ( .A(n1221), .Z(n1224) );
  IVSVTX0H U428 ( .A(n1000), .Z(n827) );
  ND3SVTX2 U429 ( .A(n1378), .B(n511), .C(n509), .Z(n1405) );
  NR2SVTX2 U430 ( .A(n1408), .B(n259), .Z(n532) );
  ND3SVTX6 U431 ( .A(n389), .B(n390), .C(n799), .Z(n539) );
  ND4ASVTX4 U432 ( .A(n1461), .B(n1462), .C(n1434), .D(n375), .Z(n493) );
  IVSVTX6 U433 ( .A(n1230), .Z(n281) );
  IVSVTX2 U434 ( .A(n1462), .Z(n263) );
  IVSVTX2 U435 ( .A(n1487), .Z(n390) );
  IVSVTX2 U436 ( .A(n1179), .Z(n460) );
  IVSVTX2 U437 ( .A(n1259), .Z(n1260) );
  NR2SVTX4 U438 ( .A(n218), .B(n791), .Z(n799) );
  CTBUFSVTX2 U439 ( .A(n1468), .Z(n348) );
  IVSVTX4 U440 ( .A(n287), .Z(n262) );
  AO4SVTX2 U441 ( .A(n1369), .B(n1466), .C(O[27]), .D(n1368), .Z(n1409) );
  F_ND2ASVTX2 U442 ( .A(n1345), .B(n1357), .Z(n1523) );
  ND3ABSVTX4 U443 ( .A(n1229), .B(n589), .C(n337), .Z(n752) );
  IVSVTX1 U444 ( .A(n1248), .Z(n216) );
  IVSVTX6 U445 ( .A(n1391), .Z(n1000) );
  ND2ASVTX6 U446 ( .A(n1496), .B(n1506), .Z(n1526) );
  ND2ASVTX6 U447 ( .A(n1367), .B(n1366), .Z(n1408) );
  IVSVTX2 U448 ( .A(n1346), .Z(n1357) );
  ND2ASVTX6 U449 ( .A(n584), .B(n1379), .Z(n821) );
  IVSVTX2 U450 ( .A(n1270), .Z(n285) );
  CTIVSVTX4 U451 ( .A(n611), .Z(n1497) );
  IVSVTX4 U452 ( .A(n1345), .Z(n1327) );
  AN2SVTX1 U453 ( .A(n412), .B(n1176), .Z(n875) );
  NR2SVTX2 U454 ( .A(n1177), .B(n1183), .Z(n1142) );
  ND2ASVTX4 U455 ( .A(n364), .B(n1326), .Z(n362) );
  IVSVTX2 U456 ( .A(n1488), .Z(n218) );
  AO7ABSVTX6 U457 ( .A(n1467), .B(n1466), .C(n1465), .Z(n1502) );
  IVSVTX6 U458 ( .A(n266), .Z(n589) );
  IVSVTX4 U459 ( .A(n1424), .Z(n290) );
  BFSVTX4 U460 ( .A(n1211), .Z(n1141) );
  ND2SVTX6 U461 ( .A(n1212), .B(n1243), .Z(n1227) );
  CTBUFSVTX2 U462 ( .A(n1332), .Z(n354) );
  NR3SVTX4 U463 ( .A(n1490), .B(n289), .C(n1499), .Z(n1485) );
  AO7SVTX4 U464 ( .A(n1427), .B(n1422), .C(n1421), .Z(n1461) );
  AO39SVTX6 U465 ( .A(n1182), .B(n309), .C(n1181), .D(n240), .E(n753), .F(
        n1180), .Z(n1251) );
  IVSVTX6 U466 ( .A(n266), .Z(n723) );
  ND2SVTX2 U467 ( .A(n1365), .B(n1477), .Z(n1481) );
  IVSVTX12 U468 ( .A(n251), .Z(n1475) );
  BFSVTX6 U469 ( .A(n1207), .Z(n240) );
  ND3ASVTX4 U470 ( .A(n1365), .B(n1472), .C(n1473), .Z(n1474) );
  F_ND2ASVTX2 U471 ( .A(n1466), .B(n1464), .Z(n1465) );
  AO4SVTX2 U472 ( .A(n1183), .B(n1181), .C(n1177), .D(n1195), .Z(n975) );
  AO2SVTX4 U473 ( .A(n1198), .B(n470), .C(n412), .D(n759), .Z(n469) );
  IVSVTX2 U474 ( .A(n1473), .Z(n324) );
  IVSVTX2 U475 ( .A(n1174), .Z(n759) );
  ND2ASVTX6 U476 ( .A(n251), .B(n231), .Z(n1038) );
  ND2SVTX4 U477 ( .A(n1440), .B(n1441), .Z(n585) );
  B_IVSVTX1 U478 ( .A(n1194), .Z(n1177) );
  ND2SVTX6 U479 ( .A(O[27]), .B(n1210), .Z(n1158) );
  ND3SVTX6 U480 ( .A(n509), .B(n864), .C(n1378), .Z(n364) );
  CTIVSVTX6 U481 ( .A(n1183), .Z(n471) );
  ND3SVTX2 U482 ( .A(O[27]), .B(n1283), .C(n1282), .Z(n1285) );
  CTBUFSVTX4 U483 ( .A(n1363), .Z(n232) );
  ND2ASVTX6 U484 ( .A(n1204), .B(n1175), .Z(n1284) );
  NR2SVTX2 U485 ( .A(n1180), .B(n1207), .Z(n719) );
  IVSVTX6 U486 ( .A(n1195), .Z(n412) );
  ND2ASVTX6 U487 ( .A(n398), .B(n1168), .Z(n570) );
  F_IVSVTX1 U488 ( .A(n1184), .Z(n1174) );
  ND2SVTX2 U489 ( .A(n1176), .B(n654), .Z(n758) );
  NR2SVTX6 U490 ( .A(n215), .B(n1207), .Z(n1470) );
  ND2SVTX6 U491 ( .A(n550), .B(n549), .Z(n1432) );
  IVSVTX8 U492 ( .A(n1363), .Z(O[27]) );
  ND2SVTX2 U493 ( .A(n1175), .B(n292), .Z(n757) );
  CTIVSVTX2 U494 ( .A(n509), .Z(n676) );
  B_ND2SVTX2 U495 ( .A(n1191), .B(n230), .Z(n1172) );
  BFSVTX2 U496 ( .A(n1169), .Z(n383) );
  BFSVTX4 U497 ( .A(n1128), .Z(n215) );
  B_IVSVTX1 U498 ( .A(n1427), .Z(n230) );
  IVSVTX0H U499 ( .A(n1151), .Z(n961) );
  IVSVTX4 U500 ( .A(n1206), .Z(n269) );
  ND2SVTX2 U501 ( .A(n941), .B(n1184), .Z(n325) );
  ND2SVTX2 U502 ( .A(n1098), .B(n1099), .Z(n1126) );
  ND2SVTX4 U503 ( .A(n1091), .B(n1392), .Z(n690) );
  IVSVTX4 U504 ( .A(n1116), .Z(n735) );
  ND2SVTX6 U505 ( .A(n247), .B(n546), .Z(n548) );
  ND2SVTX4 U506 ( .A(n730), .B(n1090), .Z(n629) );
  ND2SVTX6 U507 ( .A(n724), .B(O[28]), .Z(n1330) );
  NR2ASVTX6 U508 ( .A(n251), .B(n1129), .Z(n1507) );
  IVSVTX1 U509 ( .A(n1106), .Z(n1166) );
  ND2SVTX6 U510 ( .A(n326), .B(n651), .Z(n1382) );
  AO7ABSVTX4 U511 ( .A(n1096), .B(n1095), .C(n1311), .Z(n400) );
  AO17SVTX4 U512 ( .A(n1007), .B(n1169), .C(n1147), .D(n712), .Z(n555) );
  NR2SVTX2 U513 ( .A(n941), .B(n942), .Z(n943) );
  F_IVSVTX1 U514 ( .A(n271), .Z(n724) );
  BFSVTX4 U515 ( .A(n1204), .Z(n309) );
  CTIVSVTX6 U516 ( .A(n1091), .Z(n326) );
  ND2ASVTX6 U517 ( .A(n1082), .B(n1155), .Z(n829) );
  IVSVTX6 U518 ( .A(n1450), .Z(n544) );
  IVSVTX2 U519 ( .A(n957), .Z(n347) );
  ND2SVTX4 U520 ( .A(n951), .B(n950), .Z(n1176) );
  IVSVTX0H U521 ( .A(n1150), .Z(n958) );
  CTIVSVTX2 U522 ( .A(n515), .Z(n1182) );
  IVSVTX8 U523 ( .A(n1311), .Z(n1009) );
  NR3ABSVTX6 U524 ( .A(N[0]), .B(n1119), .C(n1118), .Z(n546) );
  IVSVTX2 U525 ( .A(n1090), .Z(n651) );
  IVSVTX8 U526 ( .A(n1128), .Z(n268) );
  NR3ASVTX2 U527 ( .A(n843), .B(n941), .C(n1205), .Z(n969) );
  IVSVTX1 U528 ( .A(n1167), .Z(n558) );
  ND2ASVTX4 U529 ( .A(n271), .B(n710), .Z(n998) );
  AO20SVTX4 U530 ( .A(n1067), .B(n1077), .C(O[29]), .D(n1375), .Z(n1068) );
  CTIVSVTX2 U531 ( .A(n1322), .Z(n778) );
  CTIVSVTX2 U532 ( .A(n1070), .Z(n1082) );
  ND2ASVTX6 U533 ( .A(n273), .B(n957), .Z(n1151) );
  ND2SVTX4 U534 ( .A(n1056), .B(n1057), .Z(n1063) );
  CTIVSVTX2 U535 ( .A(n1146), .Z(n410) );
  AO7ASVTX4 U536 ( .A(n860), .B(n633), .C(n588), .Z(n1138) );
  IVSVTX4 U537 ( .A(n1096), .Z(n1375) );
  AO2SVTX2 U538 ( .A(n1106), .B(n1019), .C(n1119), .D(n1144), .Z(n939) );
  ND2SVTX2 U539 ( .A(n1103), .B(n1029), .Z(n1152) );
  ND3SVTX4 U540 ( .A(n1028), .B(n602), .C(n601), .Z(n1202) );
  NR3SVTX4 U541 ( .A(n1830), .B(n296), .C(n825), .Z(n1140) );
  ND2ASVTX4 U542 ( .A(O[29]), .B(n515), .Z(n1137) );
  F_ND2ASVTX2 U543 ( .A(n272), .B(n1121), .Z(n1122) );
  NR2ASVTX4 U544 ( .A(n1101), .B(n1830), .Z(n1150) );
  BFSVTX0H U545 ( .A(n949), .Z(n310) );
  IVSVTX2 U546 ( .A(n1119), .Z(n935) );
  IVSVTX0H U547 ( .A(n273), .Z(n848) );
  ND2SVTX2 U548 ( .A(n1025), .B(n1163), .Z(n1028) );
  AO7SVTX4 U549 ( .A(n273), .B(n673), .C(n687), .Z(n993) );
  IVSVTX4 U550 ( .A(n994), .Z(n987) );
  ND2SVTX4 U551 ( .A(n1060), .B(n1084), .Z(n1061) );
  ND2SVTX6 U552 ( .A(n997), .B(n415), .Z(n732) );
  AO7ABSVTX4 U553 ( .A(n988), .B(n1064), .C(n1058), .Z(n1062) );
  NR3ABSVTX4 U554 ( .A(n860), .B(n252), .C(n1030), .Z(n522) );
  ND2ASVTX6 U555 ( .A(n1072), .B(n1012), .Z(n1096) );
  IVSVTX4 U556 ( .A(n1136), .Z(n514) );
  AO7CSVTX6 U557 ( .A(n1097), .B(n1008), .C(n1007), .Z(n1094) );
  ND2SVTX6 U558 ( .A(n985), .B(n986), .Z(n994) );
  NR2SVTX6 U559 ( .A(n294), .B(n244), .Z(n523) );
  AO7SVTX6 U560 ( .A(n989), .B(n990), .C(n688), .Z(n997) );
  ND2ASVTX6 U561 ( .A(n630), .B(n244), .Z(n402) );
  IVSVTX10 U562 ( .A(n733), .Z(n1007) );
  ND3SVTX6 U563 ( .A(N[3]), .B(n632), .C(n1029), .Z(n1079) );
  ND3ABSVTX4 U564 ( .A(n860), .B(n1015), .C(n1030), .Z(n1066) );
  ND2SVTX2 U565 ( .A(n1161), .B(n1830), .Z(n1032) );
  AO4ABSVTX4 U566 ( .C(n825), .D(n1016), .A(N[10]), .B(n688), .Z(n401) );
  IVSVTX0H U567 ( .A(N[24]), .Z(n945) );
  ND2SVTX1 U568 ( .A(n1161), .B(n1006), .Z(n985) );
  IVSVTX0H U569 ( .A(n1027), .Z(n399) );
  BFSVTX0H U570 ( .A(N[5]), .Z(n1019) );
  AO6SVTX4 U571 ( .A(n911), .B(n609), .C(n630), .Z(n693) );
  ND3ABSVTX2 U572 ( .A(n1072), .B(n838), .C(n711), .Z(n674) );
  BFSVTX10 U573 ( .A(n944), .Z(n1830) );
  ND3ABSVTX2 U574 ( .A(n1161), .B(n298), .C(n910), .Z(n911) );
  ND4ABSVTX6 U575 ( .A(n928), .B(n1120), .C(n953), .D(n838), .Z(n694) );
  IVSVTX8 U576 ( .A(n978), .Z(n838) );
  IVSVTX6 U577 ( .A(n980), .Z(n743) );
  IVSVTX6 U578 ( .A(n983), .Z(n1006) );
  ND2SVTX6 U579 ( .A(n927), .B(n811), .Z(n706) );
  BFSVTX2 U580 ( .A(N[17]), .Z(n953) );
  AO4SVTX2 U581 ( .A(n900), .B(n909), .C(n1160), .D(n890), .Z(n610) );
  BFSVTX2 U582 ( .A(N[6]), .Z(n1161) );
  BFSVTX2 U583 ( .A(N[8]), .Z(n1025) );
  ND2SVTX6 U584 ( .A(n934), .B(n1041), .Z(n982) );
  NR3ABSVTX6 U585 ( .A(n834), .B(n738), .C(n984), .Z(n907) );
  NR2SVTX2 U586 ( .A(n295), .B(n851), .Z(n905) );
  ND2SVTX2 U587 ( .A(n1015), .B(N[9]), .Z(n909) );
  BFSVTX2 U588 ( .A(N[22]), .Z(n1162) );
  ND2ASVTX6 U589 ( .A(n949), .B(n929), .Z(n931) );
  IVSVTX2 U590 ( .A(N[6]), .Z(n1072) );
  ND3SVTX6 U591 ( .A(n894), .B(n892), .C(n893), .Z(n895) );
  IVSVTX2 U592 ( .A(N[2]), .Z(n272) );
  BFSVTX4 U593 ( .A(N[7]), .Z(n1083) );
  IVSVTX2 U594 ( .A(n1015), .Z(n524) );
  NR2SVTX6 U595 ( .A(n843), .B(n916), .Z(n314) );
  NR2SVTX6 U596 ( .A(n914), .B(n918), .Z(n934) );
  BFSVTX2 U597 ( .A(N[18]), .Z(n1120) );
  BFSVTX2 U598 ( .A(N[19]), .Z(n1103) );
  ND2SVTX4 U599 ( .A(N[11]), .B(n890), .Z(n891) );
  IVSVTX2 U600 ( .A(N[25]), .Z(n954) );
  IVSVTX4 U601 ( .A(N[26]), .Z(n949) );
  NR2SVTX6 U602 ( .A(N[20]), .B(N[21]), .Z(n1013) );
  NR2SVTX6 U603 ( .A(N[27]), .B(N[24]), .Z(n715) );
  CTBUFSVTX8 U604 ( .A(n1696), .Z(n377) );
  IVSVTX4 U605 ( .A(n377), .Z(n1697) );
  EOSVTX8 U606 ( .A(n1699), .B(n1698), .Z(O[19]) );
  AO4ABSVTX6 U607 ( .C(n1561), .D(n472), .A(n1558), .B(n861), .Z(n341) );
  NR2SVTX6 U608 ( .A(n1083), .B(n941), .Z(n1085) );
  BFSVTX4 U609 ( .A(n1513), .Z(n211) );
  IVSVTX4 U610 ( .A(n212), .Z(n1315) );
  NR2SVTX4 U611 ( .A(n1475), .B(n1313), .Z(n212) );
  CTIVSVTX4 U612 ( .A(n1047), .Z(n709) );
  IVSVTX8 U613 ( .A(n299), .Z(n1341) );
  BFSVTX10 U614 ( .A(n820), .Z(n385) );
  ND2SVTX6 U615 ( .A(n542), .B(n1469), .Z(n537) );
  NR2SVTX6 U616 ( .A(n1480), .B(n1100), .Z(n302) );
  ND2SVTX4 U617 ( .A(n1376), .B(n213), .Z(n1049) );
  NR2SVTX4 U618 ( .A(n251), .B(n1143), .Z(n213) );
  ND2ASVTX8 U619 ( .A(O[29]), .B(n823), .Z(n1143) );
  IVSVTX8 U620 ( .A(n589), .Z(n375) );
  AN2SVTX8 U621 ( .A(n266), .B(n1370), .Z(n1371) );
  IVSVTX12 U622 ( .A(n1143), .Z(n291) );
  IVSVTX10 U623 ( .A(n291), .Z(n657) );
  ND3SVTX8 U624 ( .A(n1493), .B(n660), .C(n1492), .Z(n356) );
  IVSVTX6 U625 ( .A(n356), .Z(n407) );
  IVSVTX8 U626 ( .A(n311), .Z(n1235) );
  BFSVTX8 U627 ( .A(n1030), .Z(n386) );
  ND3SVTX8 U628 ( .A(n1506), .B(n1502), .C(n214), .Z(n1503) );
  NR3SVTX6 U629 ( .A(n579), .B(n1500), .C(n1499), .Z(n214) );
  NR2SVTX6 U630 ( .A(N[26]), .B(N[25]), .Z(n714) );
  CTIVSVTX4 U631 ( .A(N[23]), .Z(n843) );
  AO7SVTX8 U632 ( .A(n1597), .B(n1304), .C(n1300), .Z(n447) );
  ND2SVTX6 U633 ( .A(n1533), .B(n796), .Z(n1716) );
  IVSVTX10 U634 ( .A(n1047), .Z(n823) );
  IVSVTX8 U635 ( .A(n978), .Z(n235) );
  IVSVTX8 U636 ( .A(n314), .Z(n868) );
  IVSVTX12 U637 ( .A(n726), .Z(n686) );
  AO2SVTX8 U638 ( .A(n728), .B(n1059), .C(n686), .D(n993), .Z(n1392) );
  AO7SVTX6 U639 ( .A(n988), .B(n689), .C(n981), .Z(n1059) );
  NR2ASVTX6 U640 ( .A(n216), .B(n1269), .Z(n1275) );
  NR3SVTX8 U641 ( .A(n1266), .B(n367), .C(n1248), .Z(n816) );
  IVSVTX8 U642 ( .A(n1256), .Z(n646) );
  AO7CSVTX6 U643 ( .A(n257), .B(n646), .C(n1228), .Z(n665) );
  AO4SVTX4 U644 ( .A(n1285), .B(n1186), .C(n1475), .D(n1480), .Z(n1286) );
  IVSVTX8 U645 ( .A(n952), .Z(n1207) );
  AN2SVTX8 U646 ( .A(n1063), .B(n952), .Z(n1321) );
  AO2ABSVTX8 U647 ( .C(n385), .D(n1494), .A(n1823), .B(n1493), .Z(n465) );
  ND3SVTX8 U648 ( .A(n1363), .B(n1063), .C(n291), .Z(n1050) );
  ND2SVTX8 U649 ( .A(n992), .B(n991), .Z(n1391) );
  IVSVTX2 U650 ( .A(n656), .Z(n1287) );
  ND2ASVTX8 U651 ( .A(n220), .B(n291), .Z(n656) );
  ND2SVTX4 U652 ( .A(n1363), .B(n268), .Z(n220) );
  NR3ABSVTX8 U653 ( .A(n1219), .B(n1173), .C(n1550), .Z(n311) );
  AO4SVTX6 U654 ( .A(n718), .B(n1365), .C(n1222), .D(n1475), .Z(n1219) );
  AO7CSVTX4 U655 ( .A(n338), .B(n1627), .C(n1626), .Z(n477) );
  ND2SVTX4 U656 ( .A(n221), .B(n1236), .Z(n1238) );
  NR2SVTX4 U657 ( .A(n1256), .B(n1235), .Z(n221) );
  IVSVTX10 U658 ( .A(n823), .Z(n712) );
  IVSVTX10 U659 ( .A(n712), .Z(n775) );
  ND3SVTX8 U660 ( .A(n1434), .B(n337), .C(n494), .Z(n1288) );
  IVSVTX4 U661 ( .A(n978), .Z(n605) );
  AN3SVTX6 U662 ( .A(n1082), .B(n1078), .C(n1079), .Z(n1087) );
  IVSVTX10 U663 ( .A(n360), .Z(n861) );
  ND2SVTX6 U664 ( .A(n1636), .B(n1629), .Z(n1630) );
  ND2ASVTX8 U665 ( .A(n823), .B(n1076), .Z(n1089) );
  ND2SVTX4 U666 ( .A(n1217), .B(n222), .Z(n1247) );
  AO7SVTX6 U667 ( .A(n223), .B(n861), .C(n432), .Z(n1611) );
  AO7ASVTX4 U668 ( .A(n266), .B(n359), .C(n263), .Z(n492) );
  AO7SVTX4 U669 ( .A(n946), .B(n1830), .C(n945), .Z(n227) );
  IVSVTX8 U670 ( .A(n1228), .Z(n248) );
  ND2ASVTX8 U671 ( .A(n1228), .B(n1510), .Z(n1527) );
  NR2SVTX6 U672 ( .A(n1650), .B(n1587), .Z(n1652) );
  IVSVTX12 U673 ( .A(n647), .Z(n929) );
  IVSVTX4 U674 ( .A(n832), .Z(n318) );
  NR2ASVTX6 U675 ( .A(n1475), .B(n1284), .Z(n1113) );
  BFSVTX1 U676 ( .A(n247), .Z(n225) );
  ND3ASVTX6 U677 ( .A(n227), .B(n948), .C(n514), .Z(n515) );
  AO2ABSVTX8 U678 ( .C(n1665), .D(n1443), .A(n263), .B(n771), .Z(n773) );
  BFSVTX1 U679 ( .A(n1804), .Z(n228) );
  IVSVTX4 U680 ( .A(n414), .Z(n1329) );
  BFSVTX10 U681 ( .A(n251), .Z(n1365) );
  IVSVTX8 U682 ( .A(n1526), .Z(n1518) );
  ND2ASVTX8 U683 ( .A(n608), .B(n1227), .Z(n1213) );
  IVSVTX10 U684 ( .A(n720), .Z(n1498) );
  IVSVTX8 U685 ( .A(n371), .Z(n952) );
  IVSVTX6 U686 ( .A(n1307), .Z(n231) );
  ND2SVTX8 U687 ( .A(n1042), .B(n1041), .Z(n944) );
  CTIVSVTX6 U688 ( .A(n1321), .Z(n1046) );
  NR2SVTX6 U689 ( .A(N[11]), .B(N[10]), .Z(n649) );
  AO20SVTX8 U690 ( .A(n234), .B(n233), .C(n1516), .D(n1234), .Z(n1245) );
  IVSVTX4 U691 ( .A(n801), .Z(n233) );
  ND2SVTX4 U692 ( .A(n1255), .B(n1236), .Z(n234) );
  IVSVTX4 U693 ( .A(n970), .Z(n971) );
  AO4SVTX6 U694 ( .A(n971), .B(n972), .C(n753), .D(n973), .Z(n744) );
  NR2SVTX4 U695 ( .A(n1010), .B(n1011), .Z(n689) );
  NR2ASVTX6 U696 ( .A(N[0]), .B(n1043), .Z(n1011) );
  IVSVTX12 U697 ( .A(n630), .Z(n860) );
  AO7SVTX6 U698 ( .A(n917), .B(n739), .C(n929), .Z(n980) );
  NR3SVTX8 U699 ( .A(n1227), .B(n489), .C(n1626), .Z(n303) );
  AO6SVTX8 U700 ( .A(n1435), .B(n248), .C(n303), .Z(n553) );
  ND3ABSVTX6 U701 ( .A(n296), .B(n838), .C(n742), .Z(n996) );
  ENSVTX8 U702 ( .A(n489), .B(n299), .Z(n1435) );
  IVSVTX8 U703 ( .A(n585), .Z(n1379) );
  ND2ASVTX8 U704 ( .A(n1450), .B(n236), .Z(n327) );
  ND2SVTX4 U705 ( .A(n1426), .B(n1004), .Z(n236) );
  ND2ASVTX8 U706 ( .A(n751), .B(n590), .Z(n1437) );
  ND3SVTX8 U707 ( .A(n237), .B(n644), .C(n643), .Z(n526) );
  BFSVTX1 U708 ( .A(n1759), .Z(n238) );
  AO1CSVTX6 U709 ( .A(n1299), .B(n594), .C(n239), .D(n372), .Z(n593) );
  IVSVTX8 U710 ( .A(n686), .Z(n728) );
  NR2SVTX4 U711 ( .A(n1453), .B(n1447), .Z(n473) );
  NR2SVTX4 U712 ( .A(n1450), .B(n1004), .Z(n1453) );
  IVSVTX10 U713 ( .A(n1621), .Z(n441) );
  IVSVTX12 U714 ( .A(n441), .Z(n446) );
  AO2SVTX8 U715 ( .A(n251), .B(n1362), .C(n612), .D(O[28]), .Z(n615) );
  ND4SVTX8 U716 ( .A(n1271), .B(n1273), .C(n1272), .D(n1274), .Z(n767) );
  IVSVTX8 U717 ( .A(n321), .Z(n791) );
  AO2SVTX8 U718 ( .A(n1178), .B(n1199), .C(n1194), .D(n654), .Z(n1187) );
  IVSVTX6 U719 ( .A(n723), .Z(n494) );
  ND3SVTX8 U720 ( .A(n469), .B(n438), .C(n436), .Z(n1291) );
  AO7ABSVTX8 U721 ( .A(n412), .B(n1197), .C(n1200), .Z(n1248) );
  ND3SVTX4 U722 ( .A(N[3]), .B(n1006), .C(n1065), .Z(n536) );
  AO7SVTX4 U723 ( .A(n1427), .B(n1426), .C(n536), .Z(n414) );
  AN2SVTX4 U724 ( .A(n412), .B(n1199), .Z(n1261) );
  ND3SVTX4 U725 ( .A(n1064), .B(n1056), .C(n1057), .Z(n1058) );
  F_ND2ASVTX2 U726 ( .A(n297), .B(n1106), .Z(n1115) );
  ND2SVTX2 U727 ( .A(N[25]), .B(n949), .Z(n582) );
  IVSVTX0H U728 ( .A(n1592), .Z(n790) );
  AO17SVTX2 U729 ( .A(O[29]), .B(n1376), .C(n1375), .D(n1428), .Z(n511) );
  IVSVTX2 U730 ( .A(n1420), .Z(n1422) );
  IVSVTX2 U731 ( .A(n1484), .Z(n1490) );
  ENSVTX1 U732 ( .A(n804), .B(n1556), .Z(n1558) );
  IVSVTX0H U733 ( .A(n1743), .Z(n1745) );
  F_ND2SVTX0H U734 ( .A(n1716), .B(n1717), .Z(n1720) );
  F_AN2SVTX2 U735 ( .A(n1601), .B(n274), .Z(n242) );
  AO6NSVTX4 U736 ( .A(n1190), .B(n1189), .C(n1466), .Z(n243) );
  IVSVTX4 U737 ( .A(n890), .Z(n841) );
  CTBUFSVTX8 U738 ( .A(N[12]), .Z(n936) );
  IVSVTX4 U739 ( .A(n1823), .Z(n379) );
  IVSVTX4 U740 ( .A(n1267), .Z(n1276) );
  IVSVTX10 U741 ( .A(n604), .Z(n978) );
  ND3ABSVTX2 U742 ( .A(n838), .B(n296), .C(n850), .Z(n981) );
  IVSVTX8 U743 ( .A(n860), .Z(n632) );
  IVSVTX12 U744 ( .A(n1029), .Z(n1030) );
  IVSVTX10 U745 ( .A(n1029), .Z(n825) );
  IVSVTX12 U746 ( .A(n402), .Z(n1106) );
  IVSVTX10 U747 ( .A(n1516), .Z(n483) );
  IVSVTX8 U748 ( .A(n483), .Z(n745) );
  IVSVTX2 U749 ( .A(n1406), .Z(n1401) );
  ND4ASVTX4 U750 ( .A(N[17]), .B(n588), .C(n959), .D(n897), .Z(n599) );
  AO2ABSVTX4 U751 ( .C(n385), .D(n1505), .A(n278), .B(n1823), .Z(n541) );
  AO2SVTX2 U752 ( .A(n1119), .B(n1134), .C(n936), .D(n1163), .Z(n938) );
  AO2SVTX4 U753 ( .A(n1119), .B(n1162), .C(n1163), .D(n1160), .Z(n950) );
  IVSVTX12 U754 ( .A(n849), .Z(n1041) );
  IVSVTX4 U755 ( .A(n726), .Z(n528) );
  ND2SVTX2 U756 ( .A(n1733), .B(n1734), .Z(n1741) );
  AO7SVTX4 U757 ( .A(n920), .B(n844), .C(n923), .Z(n456) );
  AO6SVTX4 U758 ( .A(n923), .B(n524), .C(n1160), .Z(n924) );
  NR2SVTX2 U759 ( .A(n582), .B(n647), .Z(n908) );
  NR2SVTX2 U760 ( .A(n270), .B(n1143), .Z(n1203) );
  ND3ABSVTX6 U761 ( .A(n585), .B(n584), .C(n1370), .Z(n611) );
  IVSVTX8 U762 ( .A(n1709), .Z(n559) );
  ND3ABSVTX4 U763 ( .A(n290), .B(n837), .C(n1425), .Z(n535) );
  F_ND2SVTX0H U764 ( .A(n1710), .B(n1709), .Z(n1715) );
  ND2ASVTX8 U765 ( .A(n978), .B(n915), .Z(n244) );
  IVSVTX8 U766 ( .A(N[13]), .Z(n890) );
  NR3SVTX6 U767 ( .A(n1295), .B(n1278), .C(n428), .Z(n427) );
  IVSVTX8 U768 ( .A(n944), .Z(n811) );
  IVSVTX4 U769 ( .A(n879), .Z(n880) );
  IVSVTX6 U770 ( .A(n750), .Z(n901) );
  AO7SVTX8 U771 ( .A(n276), .B(n407), .C(n459), .Z(n466) );
  NR2SVTX2 U772 ( .A(n1355), .B(n720), .Z(n1352) );
  ND3ABSVTX6 U773 ( .A(N[18]), .B(N[30]), .C(n954), .Z(n919) );
  IVSVTX12 U774 ( .A(n251), .Z(n247) );
  IVSVTX6 U775 ( .A(n613), .Z(n612) );
  IVSVTX12 U776 ( .A(n451), .Z(n660) );
  AO7ABSVTX8 U777 ( .A(n1357), .B(n1327), .C(n1356), .Z(n1358) );
  AO6SVTX6 U778 ( .A(n1675), .B(n1658), .C(n1657), .Z(n1659) );
  AO6SVTX6 U779 ( .A(n1644), .B(n1692), .C(n1643), .Z(n1660) );
  ND4SVTX6 U780 ( .A(n1357), .B(n1371), .C(n1353), .D(n1352), .Z(n1359) );
  IVSVTX4 U781 ( .A(n703), .Z(n551) );
  AO21SVTX6 U782 ( .A(N[30]), .B(N[29]), .C(n587), .D(n896), .Z(n879) );
  IVSVTX4 U783 ( .A(N[29]), .Z(n295) );
  ND4SVTX8 U784 ( .A(n1131), .B(n1464), .C(n867), .D(n655), .Z(n1132) );
  ND3SVTX8 U785 ( .A(n1467), .B(n1117), .C(n302), .Z(n1133) );
  IVSVTX4 U786 ( .A(n1692), .Z(n1699) );
  IVSVTX2 U787 ( .A(n446), .Z(n1606) );
  ENSVTX4 U788 ( .A(n1751), .B(n1750), .Z(O[10]) );
  EOSVTX4 U789 ( .A(n1794), .B(n1793), .Z(O[4]) );
  ND2SVTX2 U790 ( .A(n1772), .B(n1756), .Z(n1761) );
  IVSVTX2 U791 ( .A(n1535), .Z(n1495) );
  ND2ASVTX4 U792 ( .A(n1228), .B(n1438), .Z(n534) );
  IVSVTX6 U793 ( .A(n258), .Z(n761) );
  ENSVTX4 U794 ( .A(n262), .B(n729), .Z(n828) );
  IVSVTX4 U795 ( .A(n1550), .Z(n257) );
  IVSVTX2 U796 ( .A(n1456), .Z(n261) );
  IVSVTX2 U797 ( .A(n1249), .Z(n1250) );
  ND3SVTX4 U798 ( .A(n1197), .B(n1466), .C(n458), .Z(n1196) );
  IVSVTX4 U799 ( .A(n1461), .Z(n246) );
  ND3SVTX4 U800 ( .A(n1126), .B(n251), .C(n291), .Z(n1484) );
  B_ND2SVTX2 U801 ( .A(n1466), .B(n1362), .Z(n1364) );
  ND2SVTX6 U802 ( .A(n938), .B(n937), .Z(n1175) );
  ND2SVTX6 U803 ( .A(n940), .B(n939), .Z(n1194) );
  IVSVTX4 U804 ( .A(n1006), .Z(n711) );
  IVSVTX4 U805 ( .A(n1120), .Z(n294) );
  IVSVTX4 U806 ( .A(n1708), .Z(n1613) );
  IVSVTX2 U807 ( .A(n442), .Z(n422) );
  IVSVTX4 U808 ( .A(n803), .Z(n1551) );
  IVSVTX6 U809 ( .A(n1758), .Z(n1793) );
  FAS1SVTX2 U810 ( .A(n1617), .B(n254), .CI(n853), .CO(n1579), .Z(n1638) );
  BFSVTX4 U811 ( .A(n1728), .Z(n370) );
  BFSVTX2 U812 ( .A(n1597), .Z(n1753) );
  ND2ASVTX4 U813 ( .A(n263), .B(n1463), .Z(n1814) );
  IVSVTX4 U814 ( .A(n245), .Z(n621) );
  IVSVTX2 U815 ( .A(n1823), .Z(n620) );
  ND2ASVTX4 U816 ( .A(n262), .B(n379), .Z(n488) );
  IVSVTX4 U817 ( .A(n1518), .Z(n781) );
  AN2SVTX4 U818 ( .A(n1224), .B(n1223), .Z(n1280) );
  ND2SVTX6 U819 ( .A(n774), .B(n1348), .Z(n1326) );
  MUX21NSVTX4 U820 ( .A(n1141), .B(n744), .S(n1365), .Z(n307) );
  IVSVTX2 U821 ( .A(n1405), .Z(n288) );
  AO4SVTX4 U822 ( .A(n874), .B(n1365), .C(n354), .D(O[27]), .Z(n533) );
  IVSVTX2 U823 ( .A(n1261), .Z(n1263) );
  IVSVTX4 U824 ( .A(n1368), .Z(n250) );
  CTIVSVTX2 U825 ( .A(n584), .Z(n863) );
  ND2SVTX4 U826 ( .A(n1363), .B(n999), .Z(n550) );
  NR2SVTX6 U827 ( .A(n878), .B(n1071), .Z(n1367) );
  ND3ABSVTX4 U828 ( .A(n711), .B(n273), .C(n710), .Z(n999) );
  IVSVTX12 U829 ( .A(n1157), .Z(n251) );
  IVSVTX4 U830 ( .A(n1202), .Z(n270) );
  ND2ASVTX4 U831 ( .A(n1072), .B(n1106), .Z(n951) );
  IVSVTX8 U832 ( .A(n506), .Z(n1128) );
  F_ND2ASVTX2 U833 ( .A(n296), .B(n1121), .Z(n937) );
  ND2SVTX8 U834 ( .A(n922), .B(n743), .Z(n733) );
  IVSVTX4 U835 ( .A(n738), .Z(n739) );
  ND3SVTX4 U836 ( .A(n831), .B(n272), .C(n920), .Z(n423) );
  IVSVTX6 U837 ( .A(n808), .Z(n920) );
  IVSVTX4 U838 ( .A(n916), .Z(n738) );
  IVSVTX4 U839 ( .A(N[16]), .Z(n898) );
  IVSVTX4 U840 ( .A(N[17]), .Z(n1110) );
  BFSVTX2 U841 ( .A(N[16]), .Z(n1027) );
  IVSVTX2 U842 ( .A(n272), .Z(n252) );
  AO7SVTX4 U843 ( .A(n377), .B(n1699), .C(n854), .Z(n1694) );
  B_ND2SVTX2 U844 ( .A(n1702), .B(n1701), .Z(n1703) );
  IVSVTX2 U845 ( .A(n1700), .Z(n1701) );
  NR2SVTX6 U846 ( .A(n1614), .B(n1615), .Z(n1700) );
  ND2SVTX4 U847 ( .A(n274), .B(n1666), .Z(n1824) );
  B_ND2SVTX2 U848 ( .A(n1244), .B(n1667), .Z(n1669) );
  IVSVTX2 U849 ( .A(n476), .Z(n475) );
  NR2ASVTX4 U850 ( .A(n1625), .B(n274), .Z(n476) );
  AO7ABSVTX2 U851 ( .A(n809), .B(n790), .C(n1591), .Z(n1593) );
  IVSVTX2 U852 ( .A(n421), .Z(n872) );
  AO7ABSVTX2 U853 ( .A(n809), .B(n1620), .C(n1606), .Z(n1608) );
  AO7ASVTX2 U854 ( .A(n1257), .B(n1606), .C(n229), .Z(n1590) );
  ENSVTX4 U855 ( .A(n1766), .B(n1765), .Z(O[5]) );
  IVSVTX6 U856 ( .A(n329), .Z(n1750) );
  ENSVTX4 U857 ( .A(n1791), .B(n1790), .Z(O[6]) );
  ENSVTX4 U858 ( .A(n1761), .B(n1760), .Z(O[8]) );
  ENSVTX4 U859 ( .A(n1777), .B(n1776), .Z(O[9]) );
  ENSVTX4 U860 ( .A(n1786), .B(n1785), .Z(O[7]) );
  NR2SVTX2 U861 ( .A(n1725), .B(n370), .Z(n1730) );
  B_ND2SVTX2 U862 ( .A(n1619), .B(n1618), .Z(n1623) );
  B_ND2SVTX2 U863 ( .A(n1723), .B(n1722), .Z(n1732) );
  EOSVTX4 U864 ( .A(n1820), .B(n1819), .Z(O[3]) );
  IVSVTX1 U865 ( .A(n495), .Z(n1744) );
  HA1SVTX4 U866 ( .A(n276), .B(n241), .CO(n1617), .S(n1635) );
  NR3ABSVTX6 U867 ( .A(n1767), .B(n1755), .C(n1759), .Z(n788) );
  ND2ASVTX6 U868 ( .A(n1240), .B(n1239), .Z(n1241) );
  B_ND2SVTX2 U869 ( .A(n606), .B(n1764), .Z(n1794) );
  B_ND2SVTX2 U870 ( .A(n1814), .B(n1796), .Z(n1799) );
  CTIVSVTX2 U871 ( .A(n228), .Z(n1805) );
  ND2SVTX6 U872 ( .A(n1419), .B(n1787), .Z(n1759) );
  AO5SVTX2 U873 ( .A(n562), .B(n1455), .C(n563), .Z(n561) );
  ND2SVTX6 U874 ( .A(n540), .B(n539), .Z(n1505) );
  B_ND2SVTX2 U875 ( .A(n483), .B(n279), .Z(n1568) );
  AO8DSVTX4 U876 ( .A(n1452), .B(n564), .C(n1451), .D(n1002), .Z(n563) );
  IVSVTX2 U877 ( .A(n1233), .Z(n696) );
  IVSVTX8 U878 ( .A(n450), .Z(n591) );
  IVSVTX6 U879 ( .A(n1516), .Z(n253) );
  CTBUFSVTX8 U880 ( .A(n1295), .Z(n450) );
  IVSVTX4 U881 ( .A(n1297), .Z(n254) );
  CTBUFSVTX8 U882 ( .A(n1228), .Z(n258) );
  IVSVTX4 U883 ( .A(n1400), .Z(n259) );
  ND3SVTX6 U884 ( .A(n1212), .B(n1159), .C(n1158), .Z(n405) );
  ND2SVTX4 U885 ( .A(n1325), .B(n1324), .Z(n774) );
  IVSVTX4 U886 ( .A(n1409), .Z(n260) );
  AO7SVTX4 U887 ( .A(n1365), .B(n250), .C(n1364), .Z(n1366) );
  ND3SVTX4 U888 ( .A(n1188), .B(n1365), .C(n1187), .Z(n755) );
  ND3SVTX4 U889 ( .A(n1284), .B(n1283), .C(n1282), .Z(n439) );
  IVSVTX4 U890 ( .A(n1344), .Z(n1369) );
  IVSVTX2 U891 ( .A(n658), .Z(n1130) );
  IVSVTX4 U892 ( .A(n1459), .Z(n264) );
  ND2SVTX4 U893 ( .A(n571), .B(n570), .Z(n569) );
  IVSVTX8 U894 ( .A(n1001), .Z(n265) );
  IVSVTX8 U895 ( .A(n751), .Z(n266) );
  B_ND2SVTX2 U896 ( .A(n1429), .B(n1428), .Z(n1430) );
  IVSVTX2 U897 ( .A(n1374), .Z(n1428) );
  AO1ABSVTX4 U898 ( .A(n889), .B(n1166), .C(n1165), .D(n572), .Z(n571) );
  NR2SVTX2 U899 ( .A(n961), .B(n960), .Z(n972) );
  ND2ASVTX4 U900 ( .A(n1073), .B(n1007), .Z(n1074) );
  NR2ASVTX4 U901 ( .A(n1007), .B(n1167), .Z(n572) );
  IVSVTX8 U902 ( .A(n988), .Z(n941) );
  NR2SVTX4 U903 ( .A(n298), .B(n734), .Z(n990) );
  IVSVTX4 U904 ( .A(n1429), .Z(n271) );
  ND3ABSVTX4 U905 ( .A(n1026), .B(n605), .C(n711), .Z(n672) );
  NR2SVTX8 U906 ( .A(n979), .B(n742), .Z(n988) );
  IVSVTX6 U907 ( .A(n928), .Z(n917) );
  IVSVTX2 U908 ( .A(n1083), .Z(n968) );
  ND2SVTX6 U909 ( .A(n898), .B(n1110), .Z(n914) );
  NR2SVTX6 U910 ( .A(N[12]), .B(N[15]), .Z(n576) );
  IVSVTX2 U911 ( .A(N[0]), .Z(n1026) );
  IVSVTX2 U912 ( .A(N[31]), .Z(n896) );
  IVSVTX6 U913 ( .A(N[3]), .Z(n273) );
  AO7SVTX4 U914 ( .A(n1674), .B(n1656), .C(n1655), .Z(n1657) );
  IVSVTX1 U915 ( .A(n1704), .Z(n1706) );
  NR2SVTX6 U916 ( .A(n1645), .B(n798), .Z(n1682) );
  ND2SVTX6 U917 ( .A(n1584), .B(n1585), .Z(n462) );
  ND2SVTX4 U918 ( .A(n1614), .B(n1615), .Z(n1702) );
  OR2SVTX2 U919 ( .A(n1825), .B(n1824), .Z(n869) );
  B_ND2SVTX2 U920 ( .A(n1669), .B(n1668), .Z(n1670) );
  ND3SVTX6 U921 ( .A(n1548), .B(n426), .C(n1549), .Z(n1562) );
  IVSVTX2 U922 ( .A(n1590), .Z(n1591) );
  F_ENSVTX2 U923 ( .A(n1609), .B(n1608), .Z(n1610) );
  IVSVTX2 U924 ( .A(n486), .Z(n485) );
  EOSVTX4 U925 ( .A(n1720), .B(n1719), .Z(O[14]) );
  EOSVTX4 U926 ( .A(n1747), .B(n1746), .Z(O[12]) );
  EOSVTX4 U927 ( .A(n1732), .B(n1731), .Z(O[15]) );
  AO6SVTX2 U928 ( .A(n1730), .B(n1750), .C(n1729), .Z(n1731) );
  AO6SVTX2 U929 ( .A(n1750), .B(n1724), .C(n1726), .Z(n1719) );
  AO6SVTX2 U930 ( .A(n1750), .B(n1739), .C(n1738), .Z(n1740) );
  AO6SVTX2 U931 ( .A(n1750), .B(n1749), .C(n1713), .Z(n1714) );
  AO6SVTX2 U932 ( .A(n1750), .B(n1745), .C(n1744), .Z(n1746) );
  B_ND2SVTX2 U933 ( .A(n870), .B(n1244), .Z(n1668) );
  EOSVTX4 U934 ( .A(n1807), .B(n1806), .Z(O[1]) );
  EOSVTX2 U935 ( .A(n1799), .B(n1798), .Z(O[2]) );
  ENSVTX4 U936 ( .A(n1822), .B(n429), .Z(O[0]) );
  AO6SVTX2 U937 ( .A(n429), .B(n1818), .C(n1817), .Z(n1819) );
  BFSVTX2 U938 ( .A(n1584), .Z(n857) );
  AO6SVTX2 U939 ( .A(n429), .B(n1821), .C(n1805), .Z(n1806) );
  AO5SVTX2 U940 ( .A(n1557), .B(n802), .C(n1556), .Z(n803) );
  IVSVTX8 U941 ( .A(n328), .Z(n1540) );
  IVSVTX2 U942 ( .A(n852), .Z(n853) );
  IVSVTX4 U943 ( .A(n1545), .Z(n1301) );
  B_ND2SVTX2 U944 ( .A(n1769), .B(n1772), .Z(n1775) );
  IVSVTX1 U945 ( .A(n431), .Z(n1773) );
  B_ND2SVTX2 U946 ( .A(n1753), .B(n1599), .Z(n1754) );
  B_ND2SVTX2 U947 ( .A(n1742), .B(n396), .Z(n1747) );
  IVSVTX4 U948 ( .A(n822), .Z(n780) );
  IVSVTX2 U949 ( .A(n1797), .Z(n429) );
  CTIVSVTX2 U950 ( .A(n1752), .Z(n1599) );
  B_ND2SVTX2 U951 ( .A(n346), .B(n1787), .Z(n1784) );
  B_ND2SVTX2 U952 ( .A(n1781), .B(n346), .Z(n1791) );
  IVSVTX1 U953 ( .A(n312), .Z(n1815) );
  B_ND2SVTX2 U954 ( .A(n1821), .B(n228), .Z(n1822) );
  B_ND2SVTX2 U955 ( .A(n1810), .B(n1809), .Z(n1820) );
  ND2ASVTX6 U956 ( .A(n1557), .B(n668), .Z(n667) );
  IVSVTX4 U957 ( .A(n666), .Z(n619) );
  IVSVTX6 U958 ( .A(n516), .Z(n1764) );
  ND2SVTX6 U959 ( .A(n481), .B(n480), .Z(n1525) );
  AO7SVTX4 U960 ( .A(n1557), .B(n663), .C(n695), .Z(n662) );
  IVSVTX2 U961 ( .A(n696), .Z(n574) );
  NR2ASVTX6 U962 ( .A(n263), .B(n1463), .Z(n1795) );
  IVSVTX4 U963 ( .A(n1288), .Z(n652) );
  IVSVTX4 U964 ( .A(n1235), .Z(n1225) );
  ND2SVTX4 U965 ( .A(n1386), .B(n532), .Z(n531) );
  IVSVTX4 U966 ( .A(n1442), .Z(n1445) );
  ENSVTX6 U967 ( .A(n355), .B(n535), .Z(n1438) );
  IVSVTX2 U968 ( .A(n257), .Z(n695) );
  IVSVTX2 U969 ( .A(n1523), .Z(n1347) );
  IVSVTX8 U970 ( .A(n1213), .Z(n820) );
  IVSVTX6 U971 ( .A(n336), .Z(n337) );
  IVSVTX2 U972 ( .A(n1625), .Z(n1663) );
  IVSVTX8 U973 ( .A(n1326), .Z(n282) );
  IVSVTX4 U974 ( .A(n1524), .Z(n283) );
  NR3SVTX4 U975 ( .A(n1249), .B(n1261), .C(n1221), .Z(n1208) );
  ND2ASVTX6 U976 ( .A(n716), .B(n1198), .Z(n1200) );
  IVSVTX2 U977 ( .A(n1416), .Z(n286) );
  IVSVTX4 U978 ( .A(n265), .Z(n547) );
  IVSVTX4 U979 ( .A(n364), .Z(n1349) );
  IVSVTX6 U980 ( .A(n1350), .Z(n287) );
  ND2SVTX6 U981 ( .A(n1050), .B(n1049), .Z(n1306) );
  CTIVSVTX2 U982 ( .A(n1457), .Z(n812) );
  IVSVTX4 U983 ( .A(n1483), .Z(n289) );
  IVSVTX2 U984 ( .A(n1336), .Z(n424) );
  IVSVTX2 U985 ( .A(n1284), .Z(n1186) );
  ND2SVTX6 U986 ( .A(n943), .B(n710), .Z(n1195) );
  IVSVTX10 U987 ( .A(n1118), .Z(n292) );
  ND2SVTX6 U988 ( .A(n1312), .B(n1094), .Z(n613) );
  IVSVTX4 U989 ( .A(n308), .Z(n1376) );
  IVSVTX4 U990 ( .A(n1004), .Z(n1005) );
  IVSVTX4 U991 ( .A(n1392), .Z(n510) );
  ND2ASVTX6 U992 ( .A(n1070), .B(n737), .Z(n736) );
  IVSVTX2 U993 ( .A(n674), .Z(n1073) );
  IVSVTX4 U994 ( .A(n922), .Z(n979) );
  BFSVTX2 U995 ( .A(n1830), .Z(O[31]) );
  IVSVTX2 U996 ( .A(n836), .Z(n962) );
  IVSVTX4 U997 ( .A(n1830), .Z(n293) );
  ND4ABSVTX6 U998 ( .A(n273), .B(n921), .C(n920), .D(n899), .Z(n903) );
  IVSVTX2 U999 ( .A(n936), .Z(n633) );
  NR2SVTX6 U1000 ( .A(n600), .B(n599), .Z(n1042) );
  IVSVTX2 U1001 ( .A(N[9]), .Z(n1107) );
  NR2SVTX6 U1002 ( .A(N[14]), .B(N[13]), .Z(n575) );
  BFSVTX2 U1003 ( .A(N[21]), .Z(n1144) );
  BFSVTX2 U1004 ( .A(N[20]), .Z(n1134) );
  IVSVTX6 U1005 ( .A(N[4]), .Z(n296) );
  IVSVTX4 U1006 ( .A(N[1]), .Z(n297) );
  IVSVTX4 U1007 ( .A(N[5]), .Z(n298) );
  ND3ABSVTX8 U1008 ( .A(n837), .B(n543), .C(n1331), .Z(n299) );
  IVSVTX4 U1009 ( .A(n300), .Z(n1053) );
  ND2SVTX4 U1010 ( .A(n1318), .B(n1046), .Z(n300) );
  IVSVTX8 U1011 ( .A(n1214), .Z(n1294) );
  ND2ASVTX8 U1012 ( .A(n767), .B(n762), .Z(n350) );
  AO17SVTX6 U1013 ( .A(n1072), .B(n926), .C(n925), .D(n924), .Z(n927) );
  NR2SVTX4 U1014 ( .A(n1182), .B(n753), .Z(n793) );
  ND2SVTX4 U1015 ( .A(n1475), .B(n301), .Z(n1131) );
  ND2SVTX4 U1016 ( .A(n1283), .B(n1282), .Z(n301) );
  NR2ASVTX6 U1017 ( .A(n246), .B(n1460), .Z(n1436) );
  ND2SVTX4 U1018 ( .A(n814), .B(n1262), .Z(n367) );
  AO2SVTX6 U1019 ( .A(n1178), .B(n269), .C(n1205), .D(n654), .Z(n814) );
  ND2SVTX4 U1020 ( .A(n1101), .B(n1163), .Z(n1102) );
  ND3SVTX8 U1021 ( .A(n400), .B(n304), .C(n1017), .Z(n527) );
  ND2ASVTX8 U1022 ( .A(n1312), .B(n1009), .Z(n304) );
  ENSVTX8 U1023 ( .A(n1403), .B(n1402), .Z(n1404) );
  ND3SVTX6 U1024 ( .A(n659), .B(n658), .C(n656), .Z(n349) );
  ND2SVTX4 U1025 ( .A(n291), .B(n305), .Z(n658) );
  NR2SVTX4 U1026 ( .A(n1363), .B(n1033), .Z(n305) );
  ND3ABSVTX8 U1027 ( .A(n875), .B(n1142), .C(n307), .Z(n1244) );
  NR2SVTX4 U1028 ( .A(n589), .B(n645), .Z(n1394) );
  ND3SVTX8 U1029 ( .A(n274), .B(n701), .C(n700), .Z(n1631) );
  IVSVTX4 U1030 ( .A(n984), .Z(n983) );
  NR2SVTX4 U1031 ( .A(n1067), .B(n1077), .Z(n308) );
  CTIVSVTX6 U1032 ( .A(n728), .Z(n392) );
  NR2SVTX2 U1033 ( .A(n1312), .B(n1065), .Z(n1317) );
  NR2SVTX4 U1034 ( .A(n836), .B(n978), .Z(n963) );
  AN2SVTX8 U1035 ( .A(n1493), .B(n1276), .Z(n1274) );
  BFSVTX12 U1036 ( .A(n1363), .Z(n1466) );
  BFSVTX1 U1037 ( .A(n1813), .Z(n312) );
  ND2SVTX8 U1038 ( .A(n735), .B(n387), .Z(n1024) );
  ND2SVTX8 U1039 ( .A(n1079), .B(n1078), .Z(n1322) );
  ND2SVTX6 U1040 ( .A(n1382), .B(n323), .Z(n678) );
  ND3SVTX4 U1041 ( .A(n1096), .B(n1095), .C(n1311), .Z(n319) );
  ND2SVTX4 U1042 ( .A(n1065), .B(n1363), .Z(n1071) );
  NR4ABSVTX8 U1043 ( .A(n1516), .B(n591), .C(n747), .D(n1275), .Z(n594) );
  NR2SVTX6 U1044 ( .A(n611), .B(n720), .Z(n321) );
  AO7SVTX6 U1045 ( .A(n573), .B(n1373), .C(n1372), .Z(n682) );
  ND2ASVTX8 U1046 ( .A(n1408), .B(n680), .Z(n1755) );
  OR2SVTX2 U1047 ( .A(n1427), .B(n1426), .Z(n873) );
  IVSVTX4 U1048 ( .A(n1229), .Z(n1434) );
  ND2SVTX2 U1049 ( .A(n246), .B(n1434), .Z(n359) );
  ND2ASVTX8 U1050 ( .A(n709), .B(n1086), .Z(n826) );
  IVSVTX6 U1051 ( .A(n528), .Z(n529) );
  AO7SVTX6 U1052 ( .A(n1011), .B(n1010), .C(n988), .Z(n1312) );
  NR2SVTX6 U1053 ( .A(n505), .B(n504), .Z(n503) );
  ND2SVTX6 U1054 ( .A(n1307), .B(n659), .Z(n874) );
  ND4ABSVTX8 U1055 ( .A(n1332), .B(n527), .C(n1039), .D(n1038), .Z(n1499) );
  IVSVTX8 U1056 ( .A(n1185), .Z(n1033) );
  AO7SVTX8 U1057 ( .A(n1032), .B(n386), .C(n1031), .Z(n1185) );
  ND2SVTX4 U1058 ( .A(n1230), .B(n418), .Z(n452) );
  IVSVTX4 U1059 ( .A(n1197), .Z(n317) );
  NR2SVTX4 U1060 ( .A(n1204), .B(n317), .Z(n1479) );
  IVSVTX2 U1061 ( .A(n728), .Z(n1084) );
  IVSVTX4 U1062 ( .A(n318), .Z(n543) );
  ND2SVTX6 U1063 ( .A(n1051), .B(n408), .Z(n394) );
  ND2SVTX6 U1064 ( .A(n378), .B(n1009), .Z(n1017) );
  ND3SVTX4 U1065 ( .A(n327), .B(n548), .C(n785), .Z(n645) );
  AO2SVTX6 U1066 ( .A(n619), .B(n668), .C(n620), .D(n621), .Z(n618) );
  IVSVTX4 U1067 ( .A(n319), .Z(n865) );
  AO2SVTX8 U1068 ( .A(n1045), .B(n1091), .C(n840), .D(n1094), .Z(n1319) );
  ND2ASVTX8 U1069 ( .A(n253), .B(n721), .Z(n331) );
  IVSVTX12 U1070 ( .A(n1065), .Z(n1311) );
  IVSVTX12 U1071 ( .A(n1155), .Z(n839) );
  ND2ASVTX8 U1072 ( .A(n573), .B(n1439), .Z(n491) );
  AO6SVTX8 U1073 ( .A(n1788), .B(n1419), .C(n322), .Z(n1770) );
  AO7SVTX8 U1074 ( .A(n1781), .B(n1778), .C(n1780), .Z(n322) );
  OR2SVTX8 U1075 ( .A(n838), .B(n1006), .Z(n673) );
  AO7SVTX8 U1076 ( .A(n483), .B(n384), .C(n541), .Z(n796) );
  ND3SVTX6 U1077 ( .A(n1382), .B(n323), .C(n679), .Z(n1351) );
  ND2SVTX8 U1078 ( .A(n614), .B(n615), .Z(n323) );
  NR3SVTX8 U1079 ( .A(n1471), .B(n1470), .C(n324), .Z(n1467) );
  AO7ABSVTX4 U1080 ( .A(n1114), .B(n1115), .C(n654), .Z(n1473) );
  AO6SVTX4 U1081 ( .A(n1116), .B(n325), .C(n712), .Z(n1471) );
  IVSVTX10 U1082 ( .A(n1207), .Z(n1178) );
  IVSVTX12 U1083 ( .A(n1204), .Z(n654) );
  AO7ABSVTX8 U1084 ( .A(n1083), .B(n1163), .C(n1021), .Z(n1184) );
  ND2SVTX6 U1085 ( .A(n1055), .B(n326), .Z(n628) );
  NR2SVTX4 U1086 ( .A(n969), .B(n326), .Z(n970) );
  ND3SVTX8 U1087 ( .A(n548), .B(n785), .C(n327), .Z(n832) );
  AO7SVTX8 U1088 ( .A(n815), .B(n1770), .C(n1415), .Z(n328) );
  NR2ASVTX6 U1089 ( .A(n1540), .B(n1712), .Z(n329) );
  ND2SVTX6 U1090 ( .A(n603), .B(n1390), .Z(n583) );
  ND2SVTX4 U1091 ( .A(n331), .B(n332), .Z(n330) );
  ND3ASVTX6 U1092 ( .A(n284), .B(n331), .C(n332), .Z(n345) );
  ND2ASVTX8 U1093 ( .A(n1401), .B(n330), .Z(n1780) );
  IVSVTX4 U1094 ( .A(n345), .Z(n1778) );
  AO2ABSVTX8 U1095 ( .C(n820), .D(n1390), .A(n771), .B(n260), .Z(n332) );
  ND2SVTX6 U1096 ( .A(n1389), .B(n583), .Z(n333) );
  ND3SVTX8 U1097 ( .A(n1388), .B(n530), .C(n531), .Z(n1389) );
  ND2SVTX6 U1098 ( .A(n334), .B(n335), .Z(n1597) );
  ND3SVTX8 U1099 ( .A(n635), .B(n637), .C(n634), .Z(n335) );
  IVSVTX2 U1100 ( .A(n278), .Z(n334) );
  NR2ASVTX6 U1101 ( .A(n278), .B(n335), .Z(n1752) );
  NR3ABSVTX8 U1102 ( .A(n1423), .B(n1424), .C(n837), .Z(n449) );
  ND3ASVTX8 U1103 ( .A(n1229), .B(n449), .C(n494), .Z(n1295) );
  IVSVTX4 U1104 ( .A(n449), .Z(n336) );
  AO7ABSVTX8 U1105 ( .A(n809), .B(n789), .C(n339), .Z(n474) );
  NR2SVTX6 U1106 ( .A(n684), .B(n340), .Z(n339) );
  ND2SVTX4 U1107 ( .A(n341), .B(n1648), .Z(n1674) );
  NR2SVTX4 U1108 ( .A(n1648), .B(n341), .Z(n1672) );
  ND2SVTX8 U1109 ( .A(n343), .B(n342), .Z(n647) );
  NR2SVTX6 U1110 ( .A(N[30]), .B(N[29]), .Z(n342) );
  NR2SVTX6 U1111 ( .A(N[31]), .B(N[28]), .Z(n343) );
  ND3SVTX8 U1112 ( .A(n288), .B(n1389), .C(n583), .Z(n346) );
  IVSVTX4 U1113 ( .A(n344), .Z(n1787) );
  ND2SVTX4 U1114 ( .A(n607), .B(n526), .Z(n344) );
  AN2SVTX8 U1115 ( .A(n346), .B(n345), .Z(n1419) );
  ND2ASVTX8 U1116 ( .A(n1827), .B(n797), .Z(n1828) );
  ND3SVTX8 U1117 ( .A(n274), .B(n279), .C(n1662), .Z(n426) );
  AO7SVTX8 U1118 ( .A(n505), .B(n502), .C(n565), .Z(n501) );
  IVSVTX10 U1119 ( .A(n1213), .Z(n1665) );
  IVSVTX2 U1120 ( .A(n1665), .Z(n520) );
  AO7SVTX6 U1121 ( .A(n1072), .B(n347), .C(n1164), .Z(n1165) );
  NR2ASVTX6 U1122 ( .A(n261), .B(n567), .Z(n504) );
  F_ND3SVTX2 U1123 ( .A(n1019), .B(n293), .C(n1029), .Z(n409) );
  ND3ABSVTX8 U1124 ( .A(n889), .B(n293), .C(n825), .Z(n1031) );
  NR2SVTX8 U1125 ( .A(n1503), .B(n1514), .Z(n1504) );
  NR2ASVTX8 U1126 ( .A(n489), .B(n487), .Z(n1808) );
  NR2SVTX4 U1127 ( .A(n349), .B(n1496), .Z(n655) );
  ND2SVTX4 U1128 ( .A(n1202), .B(n654), .Z(n659) );
  ND2ASVTX8 U1129 ( .A(n395), .B(n446), .Z(n413) );
  AO7ABSVTX4 U1130 ( .A(n292), .B(n1194), .C(n1193), .Z(n1249) );
  AO2SVTX4 U1131 ( .A(n1178), .B(n1194), .C(n383), .D(n654), .Z(n1190) );
  AO2ABSVTX8 U1132 ( .C(n350), .D(n351), .A(n1275), .B(n833), .Z(n597) );
  AO20SVTX8 U1133 ( .A(n1296), .B(n581), .C(n280), .D(n258), .Z(n351) );
  IVSVTX12 U1134 ( .A(n1065), .Z(n1155) );
  ENSVTX4 U1135 ( .A(n1552), .B(n1667), .Z(n1553) );
  AO6SVTX6 U1136 ( .A(n1621), .B(n1541), .C(n443), .Z(n1543) );
  AO7ASVTX4 U1137 ( .A(n1559), .B(n1664), .C(n1560), .Z(n1566) );
  ND2ASVTX8 U1138 ( .A(n513), .B(n512), .Z(n1378) );
  NR4ABSVTX8 U1139 ( .A(n1433), .B(n1432), .C(n547), .D(n832), .Z(n1370) );
  ND2ASVTX8 U1140 ( .A(n261), .B(n567), .Z(n502) );
  ND2ASVTX8 U1141 ( .A(n1213), .B(n819), .Z(n463) );
  ENSVTX8 U1142 ( .A(n283), .B(n353), .Z(n1512) );
  ND4SVTX8 U1143 ( .A(n1340), .B(n1343), .C(n1342), .D(n1341), .Z(n353) );
  NR2SVTX8 U1144 ( .A(n1048), .B(n1317), .Z(n408) );
  NR2ASVTX6 U1145 ( .A(n246), .B(n1460), .Z(n1800) );
  ND3SVTX6 U1146 ( .A(n1123), .B(n1122), .C(n1124), .Z(n1197) );
  BFSVTX1 U1147 ( .A(n1423), .Z(n355) );
  ND2SVTX4 U1148 ( .A(n467), .B(n440), .Z(n1282) );
  ND2SVTX4 U1149 ( .A(n1311), .B(n357), .Z(n692) );
  ND2SVTX4 U1150 ( .A(n732), .B(n731), .Z(n357) );
  ND3SVTX8 U1151 ( .A(n1412), .B(n1411), .C(n1413), .Z(n365) );
  ND3SVTX8 U1152 ( .A(n761), .B(n670), .C(n358), .Z(n617) );
  IVSVTX8 U1153 ( .A(n717), .Z(n1118) );
  IVSVTX6 U1154 ( .A(n1291), .Z(n1493) );
  ND3ASVTX6 U1155 ( .A(N[16]), .B(n295), .C(n631), .Z(n600) );
  ND2SVTX4 U1156 ( .A(n274), .B(n1662), .Z(n360) );
  ND2SVTX4 U1157 ( .A(n1066), .B(n361), .Z(n1044) );
  IVSVTX4 U1158 ( .A(n1077), .Z(n361) );
  NR3ABSVTX8 U1159 ( .A(n252), .B(n632), .C(n825), .Z(n1077) );
  NR3ABSVTX8 U1160 ( .A(n1328), .B(n1327), .C(n362), .Z(n1342) );
  ND3SVTX8 U1161 ( .A(n1277), .B(n1276), .C(n363), .Z(n1256) );
  IVSVTX4 U1162 ( .A(n1278), .Z(n363) );
  ND2SVTX8 U1163 ( .A(n1041), .B(n1042), .Z(n630) );
  ND2SVTX6 U1164 ( .A(n1535), .B(n1534), .Z(n1722) );
  ND4ABSVTX6 U1165 ( .A(n1491), .B(n1604), .C(n1492), .D(n660), .Z(n459) );
  IVSVTX8 U1166 ( .A(n1066), .Z(n1067) );
  IVSVTX8 U1167 ( .A(n1099), .Z(n1008) );
  IVSVTX12 U1168 ( .A(n1627), .Z(n1662) );
  ND2ASVTX8 U1169 ( .A(n272), .B(n1012), .Z(n986) );
  ND2ASVTX8 U1170 ( .A(n260), .B(n365), .Z(n1768) );
  IVSVTX4 U1171 ( .A(n1486), .Z(n389) );
  ND2ASVTX8 U1172 ( .A(n366), .B(n754), .Z(n592) );
  AO7SVTX8 U1173 ( .A(n1700), .B(n434), .C(n1702), .Z(n1692) );
  AO7SVTX6 U1174 ( .A(O[27]), .B(n1334), .C(n1333), .Z(n1346) );
  BFSVTX6 U1175 ( .A(n856), .Z(n368) );
  ND2SVTX8 U1176 ( .A(n1639), .B(n1640), .Z(n1693) );
  AO7ABSVTX8 U1177 ( .A(n1003), .B(n1420), .C(n1421), .Z(n1001) );
  NR2SVTX4 U1178 ( .A(n281), .B(n1288), .Z(n859) );
  ND2SVTX4 U1179 ( .A(n1007), .B(n1047), .Z(n371) );
  IVSVTX4 U1180 ( .A(n498), .Z(n496) );
  ND3SVTX6 U1181 ( .A(n374), .B(n534), .C(n373), .Z(n1463) );
  ND2SVTX4 U1182 ( .A(n1516), .B(n828), .Z(n373) );
  ND3SVTX6 U1183 ( .A(n740), .B(n590), .C(n375), .Z(n729) );
  NR2SVTX6 U1184 ( .A(n1682), .B(n1679), .Z(n1676) );
  ND2SVTX4 U1185 ( .A(n777), .B(n1063), .Z(n1335) );
  NR3SVTX8 U1186 ( .A(n1338), .B(n1316), .C(n1319), .Z(n1054) );
  NR3SVTX8 U1187 ( .A(n251), .B(n1335), .C(n1091), .Z(n1316) );
  IVSVTX2 U1188 ( .A(n608), .Z(n1231) );
  ND2ASVTX8 U1189 ( .A(n608), .B(n404), .Z(n573) );
  IVSVTX4 U1190 ( .A(n1047), .Z(n710) );
  AO4SVTX8 U1191 ( .A(n685), .B(n748), .C(n1619), .D(n1546), .Z(n684) );
  IVSVTX4 U1192 ( .A(n1094), .Z(n378) );
  IVSVTX10 U1193 ( .A(n1244), .Z(n1237) );
  NR4ABCSVTX6 U1194 ( .A(n381), .B(n380), .C(n310), .D(n522), .Z(n1167) );
  IVSVTX4 U1195 ( .A(n523), .Z(n380) );
  ND2SVTX4 U1196 ( .A(n524), .B(n860), .Z(n381) );
  ND2SVTX6 U1197 ( .A(n1642), .B(n1641), .Z(n1690) );
  IVSVTX4 U1198 ( .A(n1494), .Z(n384) );
  IVSVTX4 U1199 ( .A(n1074), .Z(n1075) );
  NR2SVTX6 U1200 ( .A(n394), .B(n1306), .Z(n1052) );
  NR2SVTX8 U1201 ( .A(n903), .B(n902), .Z(n454) );
  NR2SVTX8 U1202 ( .A(N[26]), .B(N[31]), .Z(n631) );
  NR2SVTX8 U1203 ( .A(n1508), .B(n1514), .Z(n1509) );
  NR3SVTX8 U1204 ( .A(n835), .B(n921), .C(n919), .Z(n457) );
  BFSVTX6 U1205 ( .A(n1231), .Z(n1626) );
  ND4SVTX8 U1206 ( .A(n1330), .B(n1440), .C(n1441), .D(n1329), .Z(n751) );
  ND3ASVTX6 U1207 ( .A(n1107), .B(n1043), .C(n632), .Z(n1057) );
  CTBUFSVTX8 U1208 ( .A(n1065), .Z(n387) );
  CTBUFSVTX8 U1209 ( .A(n749), .Z(n442) );
  ND2ASVTX8 U1210 ( .A(N[28]), .B(n631), .Z(n921) );
  ND3ASVTX8 U1211 ( .A(n1507), .B(n1506), .C(n1513), .Z(n1508) );
  ND2ASVTX8 U1212 ( .A(n245), .B(n805), .Z(n1545) );
  ND2SVTX4 U1213 ( .A(n1189), .B(n1190), .Z(n1222) );
  IVSVTX10 U1214 ( .A(n1311), .Z(O[28]) );
  IVSVTX8 U1215 ( .A(n1155), .Z(n1091) );
  ND3SVTX8 U1216 ( .A(n488), .B(n491), .C(n490), .Z(n487) );
  MUX21SVTX8 U1217 ( .A(n848), .B(N[2]), .S(n686), .Z(n1420) );
  ND3ABSVTX8 U1218 ( .A(n256), .B(n769), .C(n765), .Z(n764) );
  ND3SVTX8 U1219 ( .A(n1176), .B(n232), .C(n458), .Z(n1212) );
  NR2SVTX8 U1220 ( .A(n397), .B(n1514), .Z(n1515) );
  ND3SVTX8 U1221 ( .A(n255), .B(n1618), .C(n856), .Z(n748) );
  IVSVTX4 U1222 ( .A(n1318), .Z(n1320) );
  ND4ABSVTX8 U1223 ( .A(n1355), .B(n282), .C(n1371), .D(n1498), .Z(n1356) );
  NR3SVTX8 U1224 ( .A(n1069), .B(n676), .C(n678), .Z(n675) );
  ND3SVTX8 U1225 ( .A(n268), .B(O[29]), .C(n1311), .Z(n1023) );
  IVSVTX8 U1226 ( .A(N[28]), .Z(n588) );
  IVSVTX6 U1227 ( .A(n1493), .Z(n1604) );
  ND2SVTX4 U1228 ( .A(n1197), .B(n292), .Z(n1283) );
  NR2SVTX6 U1229 ( .A(n1795), .B(n1808), .Z(n500) );
  ND3ASVTX8 U1230 ( .A(n1406), .B(n1400), .C(n1399), .Z(n1402) );
  EO3SVTX8 U1231 ( .A(n1635), .B(n1634), .C(n455), .Z(n1615) );
  IVSVTX4 U1232 ( .A(n1513), .Z(n397) );
  IVSVTX8 U1233 ( .A(n1664), .Z(n819) );
  BFSVTX1 U1234 ( .A(n703), .Z(n398) );
  NR2ASVTX8 U1235 ( .A(n888), .B(n895), .Z(n965) );
  IVSVTX4 U1236 ( .A(n1682), .Z(n1686) );
  ND2SVTX6 U1237 ( .A(n1468), .B(n1513), .Z(n451) );
  F_ND2ASVTX2 U1238 ( .A(n399), .B(n1029), .Z(n948) );
  ND2SVTX4 U1239 ( .A(n1262), .B(n1263), .Z(n1270) );
  ND2SVTX4 U1240 ( .A(n941), .B(n401), .Z(n1095) );
  ND2SVTX4 U1241 ( .A(n982), .B(n605), .Z(n1043) );
  IVSVTX6 U1242 ( .A(n749), .Z(n1571) );
  ND2SVTX6 U1243 ( .A(n1516), .B(n1519), .Z(n784) );
  ND3SVTX8 U1244 ( .A(n618), .B(n616), .C(n617), .Z(n1569) );
  ND2SVTX2 U1245 ( .A(n1492), .B(n660), .Z(n1254) );
  IVSVTX4 U1246 ( .A(n1155), .Z(n730) );
  ND3SVTX8 U1247 ( .A(n731), .B(n732), .C(n839), .Z(n1421) );
  NR2SVTX4 U1248 ( .A(n821), .B(n543), .Z(n1425) );
  ND2SVTX4 U1249 ( .A(n1813), .B(n500), .Z(n497) );
  ND2ASVTX8 U1250 ( .A(n1461), .B(n603), .Z(n568) );
  IVSVTX4 U1251 ( .A(n405), .Z(n404) );
  BFSVTX4 U1252 ( .A(n1788), .Z(n406) );
  ND3SVTX6 U1253 ( .A(n411), .B(n409), .C(n410), .Z(n1147) );
  ND2SVTX4 U1254 ( .A(n841), .B(n1106), .Z(n411) );
  IVSVTX8 U1255 ( .A(n673), .Z(n1012) );
  ND2ASVTX8 U1256 ( .A(n1107), .B(n1163), .Z(n1108) );
  IVSVTX6 U1257 ( .A(n1531), .Z(n855) );
  IVSVTX2 U1258 ( .A(n1423), .Z(n1310) );
  IVSVTX12 U1259 ( .A(n839), .Z(n840) );
  ND3ASVTX8 U1260 ( .A(n1026), .B(n247), .C(n544), .Z(n785) );
  IVSVTX8 U1261 ( .A(n1733), .Z(n1531) );
  IVSVTX8 U1262 ( .A(n829), .Z(n1048) );
  NR2SVTX4 U1263 ( .A(n281), .B(n1288), .Z(n858) );
  ND2ASVTX8 U1264 ( .A(n968), .B(n1106), .Z(n1148) );
  ND2SVTX6 U1265 ( .A(N[3]), .B(n1106), .Z(n1105) );
  IVSVTX12 U1266 ( .A(n929), .Z(n984) );
  AO3SVTX6 U1267 ( .A(n770), .B(n760), .C(n413), .D(n422), .Z(n1622) );
  IVSVTX6 U1268 ( .A(n1198), .Z(n1183) );
  ND2SVTX4 U1269 ( .A(n856), .B(n1301), .Z(n577) );
  IVSVTX4 U1270 ( .A(n725), .Z(n415) );
  ND4SVTX1 U1271 ( .A(n1152), .B(n959), .C(n941), .D(n958), .Z(n960) );
  IVSVTX4 U1272 ( .A(n417), .Z(n842) );
  ND2SVTX4 U1273 ( .A(n1056), .B(n1057), .Z(n417) );
  IVSVTX8 U1274 ( .A(n442), .Z(n685) );
  ND3SVTX8 U1275 ( .A(n1111), .B(n433), .C(n1112), .Z(n1480) );
  AO2ABSVTX8 U1276 ( .C(n1516), .D(n1281), .A(n1280), .B(n833), .Z(n595) );
  NR2ASVTX6 U1277 ( .A(n1025), .B(n838), .Z(n1010) );
  ND2SVTX4 U1278 ( .A(n1289), .B(n1297), .Z(n769) );
  IVSVTX4 U1279 ( .A(n1295), .Z(n418) );
  ND2SVTX4 U1280 ( .A(n814), .B(n1250), .Z(n1264) );
  ND2SVTX6 U1281 ( .A(n930), .B(n931), .Z(n932) );
  ND2ASVTX8 U1282 ( .A(n657), .B(n1507), .Z(n1482) );
  IVSVTX4 U1283 ( .A(n1247), .Z(n708) );
  ND3SVTX6 U1284 ( .A(n955), .B(n866), .C(n956), .Z(n1169) );
  ND2ASVTX8 U1285 ( .A(O[29]), .B(n1322), .Z(n1116) );
  NR2SVTX4 U1286 ( .A(n1296), .B(n1214), .Z(n420) );
  NR2SVTX4 U1287 ( .A(n1581), .B(n1627), .Z(n421) );
  AO7SVTX8 U1288 ( .A(n1683), .B(n1679), .C(n1680), .Z(n1675) );
  IVSVTX4 U1289 ( .A(n1254), .Z(n668) );
  AO3CDSVTX8 U1290 ( .A(n667), .B(n671), .C(n1550), .D(n483), .Z(n616) );
  NR2SVTX4 U1291 ( .A(n423), .B(n925), .Z(n913) );
  AO7SVTX8 U1292 ( .A(n1532), .B(n779), .C(n780), .Z(n1718) );
  AO7SVTX8 U1293 ( .A(n1713), .B(n559), .C(n1710), .Z(n779) );
  NR2SVTX4 U1294 ( .A(n1346), .B(n1355), .Z(n1340) );
  ND2ASVTX8 U1295 ( .A(n250), .B(n1369), .Z(n1355) );
  ND3SVTX6 U1296 ( .A(n1339), .B(n425), .C(n424), .Z(n1344) );
  NR2SVTX4 U1297 ( .A(n1337), .B(n1048), .Z(n425) );
  BFSVTX4 U1298 ( .A(n1672), .Z(n1650) );
  ENSVTX4 U1299 ( .A(n1688), .B(n1687), .Z(O[21]) );
  ND4ABCSVTX8 U1300 ( .A(n1550), .B(n1557), .C(n1256), .D(n669), .Z(n661) );
  NR2ASVTX8 U1301 ( .A(n479), .B(n1624), .Z(n1637) );
  NR2SVTX6 U1302 ( .A(n965), .B(n454), .Z(n704) );
  ND4ABSVTX8 U1303 ( .A(n281), .B(n217), .C(n427), .D(n660), .Z(n1279) );
  IVSVTX4 U1304 ( .A(n1277), .Z(n428) );
  NR2ASVTX6 U1305 ( .A(n1232), .B(n1518), .Z(n1521) );
  ND2SVTX8 U1306 ( .A(n508), .B(n1040), .Z(n800) );
  ND2ASVTX8 U1307 ( .A(n279), .B(n1662), .Z(n700) );
  ND4ABSVTX8 U1308 ( .A(n664), .B(n665), .C(n662), .D(n661), .Z(n623) );
  AO7SVTX8 U1309 ( .A(n1302), .B(n1571), .C(n577), .Z(n443) );
  BFSVTX1 U1310 ( .A(n1602), .Z(n430) );
  MUX21NSVTX8 U1311 ( .A(N[0]), .B(N[1]), .S(n529), .Z(n1004) );
  NR2ASVTX6 U1312 ( .A(n686), .B(n1075), .Z(n1076) );
  BFSVTX1 U1313 ( .A(n1770), .Z(n431) );
  ND3SVTX8 U1314 ( .A(n1371), .B(n871), .C(n1498), .Z(n795) );
  ND3ABSVTX8 U1315 ( .A(n287), .B(n677), .C(n675), .Z(n720) );
  ND2SVTX4 U1316 ( .A(n654), .B(n269), .Z(n433) );
  IVSVTX8 U1317 ( .A(n845), .Z(n923) );
  NR2SVTX4 U1318 ( .A(n835), .B(n918), .Z(n899) );
  IVSVTX4 U1319 ( .A(n435), .Z(n434) );
  F_ENSVTX2 U1320 ( .A(n435), .B(n1703), .Z(O[18]) );
  AO7SVTX6 U1321 ( .A(n1613), .B(n1704), .C(n1705), .Z(n435) );
  ENSVTX4 U1322 ( .A(n1827), .B(n797), .Z(O[25]) );
  ND2SVTX4 U1323 ( .A(n225), .B(n437), .Z(n436) );
  ND2SVTX4 U1324 ( .A(n1188), .B(n1187), .Z(n437) );
  ND2SVTX4 U1325 ( .A(n269), .B(n292), .Z(n1188) );
  ND2SVTX4 U1326 ( .A(n1466), .B(n439), .Z(n438) );
  IVSVTX4 U1327 ( .A(n468), .Z(n440) );
  AO4ABSVTX6 U1328 ( .C(n1305), .D(n648), .A(n254), .B(n1616), .Z(n445) );
  ND2ASVTX8 U1329 ( .A(n445), .B(n444), .Z(n1621) );
  ND3ABSVTX8 U1330 ( .A(n1303), .B(n1305), .C(n447), .Z(n444) );
  AO7SVTX8 U1331 ( .A(n1588), .B(n1605), .C(n1589), .Z(n749) );
  NR2SVTX8 U1332 ( .A(n1570), .B(n1302), .Z(n1541) );
  ND2SVTX8 U1333 ( .A(n1257), .B(n1258), .Z(n1570) );
  ND4ASVTX8 U1334 ( .A(n280), .B(n618), .C(n616), .D(n617), .Z(n1257) );
  IVSVTX12 U1335 ( .A(n1145), .Z(n1029) );
  IVSVTX4 U1336 ( .A(n448), .Z(n1121) );
  ND2SVTX4 U1337 ( .A(n860), .B(n244), .Z(n448) );
  ND2ASVTX8 U1338 ( .A(n978), .B(n915), .Z(n1145) );
  NR2SVTX4 U1339 ( .A(n1292), .B(n1293), .Z(n636) );
  ND2ASVTX8 U1340 ( .A(n452), .B(n660), .Z(n1293) );
  NR2SVTX4 U1341 ( .A(n963), .B(n454), .Z(n967) );
  ND2SVTX2 U1342 ( .A(n455), .B(n485), .Z(n484) );
  ND3SVTX8 U1343 ( .A(n1110), .B(n898), .C(n959), .Z(n835) );
  ND3ASVTX8 U1344 ( .A(n918), .B(n457), .C(n456), .Z(n922) );
  IVSVTX4 U1345 ( .A(n1143), .Z(n458) );
  NR2SVTX8 U1346 ( .A(n460), .B(n1260), .Z(n1491) );
  NR2SVTX6 U1347 ( .A(N[15]), .B(N[14]), .Z(n883) );
  ND2SVTX6 U1348 ( .A(n462), .B(n461), .Z(n1646) );
  AO7SVTX8 U1349 ( .A(n857), .B(n1585), .C(n1583), .Z(n461) );
  ND2SVTX8 U1350 ( .A(n463), .B(n464), .Z(n1585) );
  AO2ABSVTX6 U1351 ( .C(n1568), .D(n1664), .A(n379), .B(n274), .Z(n464) );
  AO7ABSVTX8 U1352 ( .A(n1516), .B(n466), .C(n465), .Z(n1534) );
  ND2SVTX6 U1353 ( .A(n538), .B(n537), .Z(n1494) );
  IVSVTX4 U1354 ( .A(n270), .Z(n467) );
  IVSVTX4 U1355 ( .A(n952), .Z(n468) );
  ND2ASVTX8 U1356 ( .A(n988), .B(n1047), .Z(n1204) );
  IVSVTX4 U1357 ( .A(n1033), .Z(n470) );
  NR2SVTX8 U1358 ( .A(n247), .B(n657), .Z(n1198) );
  AO2ABSVTX8 U1359 ( .C(n759), .D(n471), .A(n270), .B(n1195), .Z(n1179) );
  IVSVTX4 U1360 ( .A(n748), .Z(n1547) );
  ND3SVTX6 U1361 ( .A(n245), .B(n1246), .C(n1245), .Z(n1618) );
  AO7ASVTX8 U1362 ( .A(n1466), .B(n1210), .C(n569), .Z(n608) );
  ND3SVTX6 U1363 ( .A(n785), .B(n548), .C(n473), .Z(n1229) );
  NR2SVTX4 U1364 ( .A(n1450), .B(n1426), .Z(n1447) );
  MUX21NSVTX8 U1365 ( .A(N[2]), .B(N[1]), .S(n686), .Z(n1426) );
  ND2ASVTX8 U1366 ( .A(n983), .B(n1065), .Z(n1450) );
  ND2SVTX6 U1367 ( .A(n1537), .B(n1724), .Z(n1539) );
  NR2SVTX8 U1368 ( .A(n1743), .B(n1532), .Z(n1724) );
  EN3SVTX8 U1369 ( .A(n275), .B(n1637), .C(n1636), .Z(n1640) );
  ND3SVTX6 U1370 ( .A(n478), .B(n475), .C(n477), .Z(n1636) );
  ND2ASVTX8 U1371 ( .A(n474), .B(n1662), .Z(n1624) );
  F_ENSVTX2 U1372 ( .A(n1623), .B(n1622), .Z(n479) );
  CTIVSVTX6 U1373 ( .A(n1525), .Z(n1511) );
  AO6SVTX8 U1374 ( .A(n1510), .B(n745), .C(n482), .Z(n480) );
  NR2SVTX8 U1375 ( .A(n277), .B(n833), .Z(n482) );
  ENSVTX8 U1376 ( .A(n1535), .B(n1504), .Z(n1510) );
  ENSVTX8 U1377 ( .A(n1533), .B(n1509), .Z(n1520) );
  ND2ASVTX8 U1378 ( .A(n489), .B(n487), .Z(n1809) );
  AO7SVTX4 U1379 ( .A(n1814), .B(n1808), .C(n1809), .Z(n498) );
  IVSVTX4 U1380 ( .A(n290), .Z(n489) );
  ND2SVTX4 U1381 ( .A(n828), .B(n761), .Z(n490) );
  ND2SVTX4 U1382 ( .A(n493), .B(n492), .Z(n1443) );
  BFSVTX0H U1383 ( .A(n779), .Z(n495) );
  AO3SVTX6 U1384 ( .A(n1797), .B(n499), .C(n497), .D(n496), .Z(n1757) );
  ND2SVTX4 U1385 ( .A(n1811), .B(n500), .Z(n499) );
  NR2SVTX4 U1386 ( .A(n1436), .B(n1803), .Z(n1811) );
  NR2ASVTX6 U1387 ( .A(n264), .B(n1458), .Z(n1803) );
  AO6ASVTX8 U1388 ( .A(n561), .B(n503), .C(n501), .Z(n1797) );
  NR2ASVTX8 U1389 ( .A(n1379), .B(n566), .Z(n505) );
  ND2SVTX6 U1390 ( .A(n507), .B(n1018), .Z(n506) );
  ND3SVTX6 U1391 ( .A(n1475), .B(n268), .C(n458), .Z(n1483) );
  ND2SVTX4 U1392 ( .A(n1019), .B(n1163), .Z(n507) );
  IVSVTX4 U1393 ( .A(n811), .Z(n508) );
  ND3SVTX6 U1394 ( .A(n632), .B(n1101), .C(n1040), .Z(n1078) );
  ND2SVTX4 U1395 ( .A(n1157), .B(n1065), .Z(n1374) );
  IVSVTX4 U1396 ( .A(n1071), .Z(n512) );
  IVSVTX4 U1397 ( .A(n1092), .Z(n513) );
  AO7SVTX6 U1398 ( .A(n1007), .B(n842), .C(n1064), .Z(n1092) );
  ND2ASVTX8 U1399 ( .A(n387), .B(n510), .Z(n509) );
  ND2ASVTX8 U1400 ( .A(n253), .B(n1398), .Z(n1417) );
  ENSVTX8 U1401 ( .A(n1401), .B(n1395), .Z(n1398) );
  AO8ASVTX8 U1402 ( .A(n1397), .B(n519), .C(n1417), .D(n286), .Z(n516) );
  NR2ASVTX4 U1403 ( .A(n1405), .B(n1823), .Z(n1397) );
  AO2ABSVTX8 U1404 ( .C(n1516), .D(n1404), .A(n1823), .B(n1401), .Z(n643) );
  ND2ASVTX8 U1405 ( .A(n520), .B(n1439), .Z(n519) );
  NR2ASVTX6 U1406 ( .A(n860), .B(n1030), .Z(n957) );
  IVSVTX4 U1407 ( .A(N[14]), .Z(n889) );
  ND2ASVTX8 U1408 ( .A(n722), .B(n1522), .Z(n525) );
  IVSVTX4 U1409 ( .A(n526), .Z(n1762) );
  IVSVTX4 U1410 ( .A(n527), .Z(n1368) );
  IVSVTX4 U1411 ( .A(n726), .Z(n725) );
  AO7ABSVTX8 U1412 ( .A(n1408), .B(n1232), .C(n1387), .Z(n530) );
  ENSVTX8 U1413 ( .A(n260), .B(n791), .Z(n1390) );
  ND2SVTX4 U1414 ( .A(n533), .B(n1309), .Z(n1524) );
  ND2SVTX8 U1415 ( .A(n1231), .B(n1227), .Z(n1228) );
  ND2SVTX6 U1416 ( .A(n1330), .B(n1329), .Z(n584) );
  AO21DSVTX8 U1417 ( .A(n1486), .B(n1487), .C(n791), .D(n1488), .Z(n540) );
  IVSVTX4 U1418 ( .A(n1604), .Z(n542) );
  ND2SVTX6 U1419 ( .A(n998), .B(n247), .Z(n549) );
  ND2SVTX8 U1420 ( .A(n942), .B(n551), .Z(n1157) );
  NR2SVTX8 U1421 ( .A(n586), .B(n693), .Z(n942) );
  ND2SVTX8 U1422 ( .A(n552), .B(n553), .Z(n1460) );
  ND2SVTX4 U1423 ( .A(n812), .B(n1516), .Z(n564) );
  ND3SVTX4 U1424 ( .A(n1154), .B(n1156), .C(n1155), .Z(n554) );
  ND2SVTX8 U1425 ( .A(n555), .B(n554), .Z(n1210) );
  ND2SVTX8 U1426 ( .A(n557), .B(n556), .Z(n1211) );
  ND2ASVTX8 U1427 ( .A(n1155), .B(n1168), .Z(n556) );
  ND2SVTX4 U1428 ( .A(n558), .B(n292), .Z(n557) );
  ND2ASVTX8 U1429 ( .A(O[27]), .B(n1211), .Z(n1159) );
  ND2SVTX6 U1430 ( .A(n641), .B(n640), .Z(n560) );
  ND2ASVTX8 U1431 ( .A(n1347), .B(n560), .Z(n1709) );
  ND2SVTX6 U1432 ( .A(n784), .B(n782), .Z(n1522) );
  ND3SVTX8 U1433 ( .A(n1446), .B(n1445), .C(n1444), .Z(n566) );
  ND2SVTX6 U1434 ( .A(n568), .B(n1449), .Z(n567) );
  MUX21NSVTX8 U1435 ( .A(n1211), .B(n1210), .S(n1475), .Z(n1243) );
  ND4ABCSVTX8 U1436 ( .A(n1138), .B(n1139), .C(n1140), .D(n1137), .Z(n1168) );
  IVSVTX12 U1437 ( .A(n573), .Z(n1516) );
  ND4ABSVTX8 U1438 ( .A(n256), .B(n574), .C(n623), .D(n624), .Z(n1258) );
  IVSVTX4 U1439 ( .A(n1258), .Z(n1588) );
  IVSVTX12 U1440 ( .A(n830), .Z(n1232) );
  AO7ABSVTX8 U1441 ( .A(n1408), .B(n259), .C(n248), .Z(n1387) );
  ND4ABSVTX8 U1442 ( .A(n964), .B(n705), .C(n904), .D(n704), .Z(n703) );
  IVSVTX12 U1443 ( .A(n1157), .Z(n1363) );
  AO20SVTX8 U1444 ( .A(n933), .B(n1162), .C(n235), .D(n932), .Z(n707) );
  IVSVTX4 U1445 ( .A(n1437), .Z(n1399) );
  ND3SVTX8 U1446 ( .A(n243), .B(n1208), .C(n816), .Z(n1278) );
  ND2SVTX2 U1447 ( .A(n1456), .B(n1232), .Z(n1451) );
  ND2SVTX6 U1448 ( .A(n576), .B(n575), .Z(n845) );
  NR2SVTX4 U1449 ( .A(N[12]), .B(N[13]), .Z(n882) );
  NR2SVTX6 U1450 ( .A(N[28]), .B(N[29]), .Z(n884) );
  ND2ASVTX6 U1451 ( .A(n578), .B(n1567), .Z(n1589) );
  ND3SVTX8 U1452 ( .A(n1475), .B(n1126), .C(n458), .Z(n580) );
  ND2SVTX6 U1453 ( .A(n1483), .B(n580), .Z(n1100) );
  ND2SVTX4 U1454 ( .A(n580), .B(n1482), .Z(n579) );
  IVSVTX4 U1455 ( .A(n581), .Z(n762) );
  ND2ASVTX8 U1456 ( .A(n1295), .B(n1294), .Z(n581) );
  ND2SVTX6 U1457 ( .A(n1003), .B(n1005), .Z(n1441) );
  ND2SVTX6 U1458 ( .A(n544), .B(n1420), .Z(n1440) );
  ND2SVTX6 U1459 ( .A(n694), .B(n977), .Z(n586) );
  IVSVTX4 U1460 ( .A(N[27]), .Z(n959) );
  ND2SVTX4 U1461 ( .A(N[27]), .B(n588), .Z(n587) );
  NR2SVTX8 U1462 ( .A(n645), .B(n837), .Z(n590) );
  ND2ASVTX8 U1463 ( .A(N[29]), .B(n897), .Z(n918) );
  NR2SVTX8 U1464 ( .A(N[19]), .B(N[24]), .Z(n897) );
  ND3SVTX8 U1465 ( .A(n1468), .B(n1230), .C(n1513), .Z(n1214) );
  ND2SVTX6 U1466 ( .A(n592), .B(n593), .Z(n1602) );
  ENSVTX8 U1467 ( .A(n254), .B(n1290), .Z(n754) );
  ND2SVTX4 U1468 ( .A(n763), .B(n764), .Z(n598) );
  ND2SVTX6 U1469 ( .A(n596), .B(n595), .Z(n1616) );
  NR2ASVTX8 U1470 ( .A(n1297), .B(n1616), .Z(n1305) );
  NR2ASVTX8 U1471 ( .A(n1491), .B(n1596), .Z(n1303) );
  AO7ASVTX8 U1472 ( .A(n745), .B(n598), .C(n597), .Z(n1596) );
  ND4ABSVTX8 U1473 ( .A(N[18]), .B(N[30]), .C(n1013), .D(n881), .Z(n849) );
  IVSVTX4 U1474 ( .A(n659), .Z(n1308) );
  ND2SVTX4 U1475 ( .A(N[0]), .B(n1121), .Z(n601) );
  ND2SVTX4 U1476 ( .A(n1027), .B(n1119), .Z(n602) );
  ND2SVTX8 U1477 ( .A(n745), .B(n1512), .Z(n1413) );
  IVSVTX10 U1478 ( .A(n1040), .Z(n1163) );
  ND2SVTX8 U1479 ( .A(n982), .B(n235), .Z(n1040) );
  NR2SVTX8 U1480 ( .A(n916), .B(n647), .Z(n604) );
  NR2ASVTX4 U1481 ( .A(n830), .B(n1403), .Z(n1383) );
  ND4SVTX8 U1482 ( .A(n1158), .B(n1212), .C(n1159), .D(n608), .Z(n830) );
  NR2SVTX4 U1483 ( .A(n610), .B(n913), .Z(n609) );
  ND2SVTX6 U1484 ( .A(n1311), .B(n1092), .Z(n1362) );
  ND2SVTX6 U1485 ( .A(n1475), .B(n865), .Z(n614) );
  ND3SVTX8 U1486 ( .A(n1226), .B(n697), .C(n625), .Z(n624) );
  ND2SVTX8 U1487 ( .A(n627), .B(n626), .Z(n625) );
  IVSVTX6 U1488 ( .A(n698), .Z(n626) );
  NR2SVTX8 U1489 ( .A(n1351), .B(n1384), .Z(n1230) );
  NR2SVTX8 U1490 ( .A(n1367), .B(n1380), .Z(n679) );
  AO4SVTX8 U1491 ( .A(n1089), .B(n1088), .C(n1087), .D(n826), .Z(n1380) );
  ND2SVTX4 U1492 ( .A(n864), .B(n1378), .Z(n1069) );
  ND2SVTX6 U1493 ( .A(n1349), .B(n1350), .Z(n1384) );
  ND2SVTX8 U1494 ( .A(n629), .B(n628), .Z(n1350) );
  ND3ABSVTX8 U1495 ( .A(n860), .B(n633), .C(n1030), .Z(n1099) );
  AO6SVTX8 U1496 ( .A(n1519), .B(n248), .C(n1521), .Z(n640) );
  ENSVTX8 U1497 ( .A(n781), .B(n1515), .Z(n1519) );
  ND2SVTX8 U1498 ( .A(n745), .B(n1520), .Z(n641) );
  ND2SVTX4 U1499 ( .A(n644), .B(n643), .Z(n642) );
  AO7SVTX8 U1500 ( .A(n1764), .B(n1762), .C(n1763), .Z(n1788) );
  ND2ASVTX8 U1501 ( .A(n262), .B(n642), .Z(n1763) );
  ND3SVTX8 U1502 ( .A(n1433), .B(n1432), .C(n265), .Z(n837) );
  ND2SVTX8 U1503 ( .A(n715), .B(n714), .Z(n916) );
  NR2SVTX6 U1504 ( .A(N[8]), .B(N[9]), .Z(n650) );
  ND2SVTX6 U1505 ( .A(n650), .B(n649), .Z(n750) );
  NR4ABCSVTX6 U1506 ( .A(n1230), .B(n652), .C(n211), .D(n653), .Z(n1290) );
  ND2SVTX4 U1507 ( .A(n1289), .B(n348), .Z(n653) );
  IVSVTX4 U1508 ( .A(n1482), .Z(n1496) );
  NR3SVTX8 U1509 ( .A(n1479), .B(n1478), .C(n1476), .Z(n1464) );
  IVSVTX6 U1510 ( .A(n1255), .Z(n671) );
  IVSVTX6 U1511 ( .A(n1293), .Z(n669) );
  AO7SVTX6 U1512 ( .A(n671), .B(n1293), .C(n1557), .Z(n670) );
  NR2ASVTX6 U1513 ( .A(n1083), .B(n673), .Z(n1070) );
  ND3SVTX8 U1514 ( .A(n1423), .B(n1424), .C(n679), .Z(n677) );
  IVSVTX4 U1515 ( .A(n1407), .Z(n680) );
  ND2SVTX4 U1516 ( .A(n683), .B(n681), .Z(n1407) );
  IVSVTX4 U1517 ( .A(n682), .Z(n681) );
  ND2SVTX4 U1518 ( .A(n248), .B(n727), .Z(n683) );
  ND3ASVTX6 U1519 ( .A(n968), .B(n742), .C(n688), .Z(n687) );
  IVSVTX4 U1520 ( .A(n605), .Z(n688) );
  ND2SVTX8 U1521 ( .A(n730), .B(n1000), .Z(n1433) );
  ND2SVTX8 U1522 ( .A(n691), .B(n690), .Z(n1423) );
  ND2SVTX6 U1523 ( .A(n1391), .B(n840), .Z(n691) );
  AO7ABSVTX8 U1524 ( .A(n1009), .B(n1055), .C(n692), .Z(n1424) );
  MUX21NSVTX8 U1525 ( .A(n993), .B(n994), .S(n725), .Z(n1055) );
  NR3SVTX8 U1526 ( .A(n905), .B(n908), .C(n907), .Z(n977) );
  ND2SVTX8 U1527 ( .A(n1225), .B(n1255), .Z(n698) );
  EO3SVTX8 U1528 ( .A(n1633), .B(n1631), .C(n1632), .Z(n1641) );
  NR2SVTX4 U1529 ( .A(n699), .B(n1624), .Z(n1632) );
  AO2SVTX6 U1530 ( .A(n818), .B(n817), .C(n1577), .D(n1578), .Z(n699) );
  AO6CSVTX6 U1531 ( .A(n1627), .B(n1663), .C(n483), .Z(n701) );
  IVSVTX12 U1532 ( .A(n702), .Z(n1047) );
  NR2SVTX8 U1533 ( .A(n966), .B(n703), .Z(n702) );
  AO7SVTX8 U1534 ( .A(n868), .B(n984), .C(n880), .Z(n705) );
  NR2SVTX8 U1535 ( .A(n849), .B(n886), .Z(n964) );
  ND2SVTX8 U1536 ( .A(n706), .B(n707), .Z(n966) );
  ND2SVTX4 U1537 ( .A(n713), .B(n1547), .Z(n847) );
  IVSVTX4 U1538 ( .A(n1199), .Z(n716) );
  IVSVTX4 U1539 ( .A(n733), .Z(n734) );
  NR2SVTX8 U1540 ( .A(n1007), .B(n1047), .Z(n717) );
  MUX21NSVTX8 U1541 ( .A(n718), .B(n744), .S(n1475), .Z(n974) );
  ND2ASVTX8 U1542 ( .A(n719), .B(n792), .Z(n718) );
  ENSVTX8 U1543 ( .A(n722), .B(n795), .Z(n721) );
  ND2SVTX6 U1544 ( .A(n977), .B(n976), .Z(n726) );
  F_EOSVTX2 U1545 ( .A(n282), .B(n795), .Z(n727) );
  AN2SVTX8 U1546 ( .A(n1423), .B(n1424), .Z(n740) );
  ND2SVTX4 U1547 ( .A(n271), .B(n725), .Z(n731) );
  ND2SVTX4 U1548 ( .A(n672), .B(n996), .Z(n1429) );
  IVSVTX4 U1549 ( .A(n736), .Z(n878) );
  ND2SVTX4 U1550 ( .A(n1007), .B(n1044), .Z(n1045) );
  NR3SVTX8 U1551 ( .A(n1007), .B(n1128), .C(n1311), .Z(n1338) );
  NR2SVTX4 U1552 ( .A(n737), .B(n712), .Z(n1337) );
  ND2ASVTX8 U1553 ( .A(n1007), .B(n1322), .Z(n737) );
  NR2SVTX8 U1554 ( .A(n741), .B(n1384), .Z(n1400) );
  IVSVTX6 U1555 ( .A(n740), .Z(n741) );
  IVSVTX6 U1556 ( .A(n743), .Z(n742) );
  AO7SVTX6 U1557 ( .A(n1237), .B(n591), .C(n1516), .Z(n746) );
  IVSVTX4 U1558 ( .A(n1294), .Z(n747) );
  ND4ABSVTX8 U1559 ( .A(n750), .B(n900), .C(n1083), .D(n888), .Z(n886) );
  NR2SVTX8 U1560 ( .A(n281), .B(n752), .Z(n1492) );
  BFSVTX6 U1561 ( .A(n1118), .Z(n753) );
  ND2SVTX6 U1562 ( .A(n883), .B(n882), .Z(n900) );
  ND2SVTX4 U1563 ( .A(n1179), .B(n1259), .Z(n1267) );
  ND2SVTX4 U1564 ( .A(n756), .B(n755), .Z(n1259) );
  ND4SVTX4 U1565 ( .A(n1475), .B(n758), .C(n757), .D(n1201), .Z(n756) );
  ND2SVTX4 U1566 ( .A(n440), .B(n1197), .Z(n1201) );
  IVSVTX6 U1567 ( .A(n809), .Z(n770) );
  AO17SVTX8 U1568 ( .A(n1711), .B(n1540), .C(n1539), .D(n1538), .Z(n809) );
  AO6SVTX8 U1569 ( .A(n1718), .B(n1537), .C(n1536), .Z(n1538) );
  ND2SVTX8 U1570 ( .A(n788), .B(n1757), .Z(n1711) );
  ND2SVTX8 U1571 ( .A(n787), .B(n786), .Z(n1607) );
  ND3SVTX8 U1572 ( .A(n1275), .B(n660), .C(n1492), .Z(n766) );
  ND2ASVTX8 U1573 ( .A(n768), .B(n1274), .Z(n1296) );
  ND2SVTX4 U1574 ( .A(n285), .B(n1271), .Z(n768) );
  AO7SVTX6 U1575 ( .A(n1576), .B(n770), .C(n1575), .Z(n1577) );
  ND2SVTX6 U1576 ( .A(n772), .B(n773), .Z(n1458) );
  ND3ABSVTX8 U1577 ( .A(n777), .B(n778), .C(n775), .Z(n1051) );
  IVSVTX4 U1578 ( .A(n1125), .Z(n776) );
  ND2ASVTX8 U1579 ( .A(n777), .B(n775), .Z(n1125) );
  ND2SVTX4 U1580 ( .A(n1199), .B(n776), .Z(n1112) );
  IVSVTX4 U1581 ( .A(n941), .Z(n777) );
  AO6SVTX8 U1582 ( .A(n1512), .B(n1665), .C(n783), .Z(n782) );
  AN2BSVTX8 U1583 ( .A(n1232), .B(n283), .Z(n783) );
  NR2SVTX6 U1584 ( .A(n1752), .B(n1304), .Z(n786) );
  ENSVTX4 U1585 ( .A(n809), .B(n1754), .Z(O[16]) );
  ND2SVTX2 U1586 ( .A(n1639), .B(n1640), .Z(n854) );
  NR2SVTX4 U1587 ( .A(n794), .B(n793), .Z(n792) );
  NR2SVTX4 U1588 ( .A(n1167), .B(n309), .Z(n794) );
  NR2ASVTX6 U1589 ( .A(n277), .B(n796), .Z(n1728) );
  AO7SVTX8 U1590 ( .A(n1661), .B(n1660), .C(n1659), .Z(n797) );
  ND2SVTX6 U1591 ( .A(n1645), .B(n798), .Z(n1683) );
  ENSVTX8 U1592 ( .A(n1586), .B(n1585), .Z(n798) );
  IVSVTX12 U1593 ( .A(n800), .Z(n1119) );
  NR2ASVTX6 U1594 ( .A(n1237), .B(n1235), .Z(n801) );
  ND3SVTX8 U1595 ( .A(n1246), .B(n1241), .C(n1245), .Z(n805) );
  F_ENSVTX2 U1596 ( .A(n1557), .B(n802), .Z(n804) );
  NR2SVTX8 U1597 ( .A(n966), .B(n806), .Z(n807) );
  ND2SVTX6 U1598 ( .A(n967), .B(n976), .Z(n806) );
  IVSVTX12 U1599 ( .A(n807), .Z(n1065) );
  ND4SVTX2 U1600 ( .A(n988), .B(n843), .C(n1149), .D(n1148), .Z(n1156) );
  IVSVTX8 U1601 ( .A(n1768), .Z(n1414) );
  IVSVTX4 U1602 ( .A(n1756), .Z(n1771) );
  AO21DSVTX4 U1603 ( .A(N[14]), .B(n936), .C(n891), .D(N[15]), .Z(n893) );
  ND4ABSVTX8 U1604 ( .A(N[7]), .B(N[6]), .C(n296), .D(n298), .Z(n808) );
  AO7SVTX8 U1605 ( .A(n730), .B(n1036), .C(n1035), .Z(n1307) );
  AO7SVTX4 U1606 ( .A(n941), .B(n1034), .C(n1065), .Z(n1035) );
  AO6SVTX8 U1607 ( .A(n1692), .B(n1644), .C(n1643), .Z(n813) );
  NR2ASVTX4 U1608 ( .A(n1185), .B(n1207), .Z(n1476) );
  ENSVTX8 U1609 ( .A(n245), .B(n1279), .Z(n1281) );
  ND2SVTX4 U1610 ( .A(n1385), .B(n1383), .Z(n1388) );
  AO7SVTX2 U1611 ( .A(n1633), .B(n1632), .C(n1631), .Z(n1582) );
  ND2SVTX4 U1612 ( .A(n1767), .B(n1755), .Z(n815) );
  AO6SVTX8 U1613 ( .A(n1771), .B(n1767), .C(n1414), .Z(n1415) );
  NR2SVTX2 U1614 ( .A(n1291), .B(n1267), .Z(n1289) );
  ND4SVTX4 U1615 ( .A(n1236), .B(n1209), .C(n1225), .D(n646), .Z(n1217) );
  ND2ASVTX6 U1616 ( .A(n711), .B(n807), .Z(n1427) );
  AO7SVTX4 U1617 ( .A(n872), .B(n338), .C(n1560), .Z(n1667) );
  AO7SVTX6 U1618 ( .A(n1716), .B(n1721), .C(n1722), .Z(n1536) );
  ENSVTX8 U1619 ( .A(n1695), .B(n1694), .Z(O[20]) );
  AO7ASVTX4 U1620 ( .A(n1103), .B(n935), .C(n1102), .Z(n1104) );
  ND2SVTX4 U1621 ( .A(n1461), .B(n1460), .Z(n1801) );
  ND3SVTX8 U1622 ( .A(n1024), .B(n1023), .C(n1022), .Z(n1332) );
  IVSVTX10 U1623 ( .A(n1007), .Z(O[29]) );
  AO7ABSVTX4 U1624 ( .A(n1638), .B(n1637), .C(n1630), .Z(n1642) );
  IVSVTX4 U1625 ( .A(n1408), .Z(n1403) );
  ND3SVTX8 U1626 ( .A(n949), .B(n897), .C(n884), .Z(n885) );
  IVSVTX4 U1627 ( .A(n1577), .Z(n818) );
  IVSVTX2 U1628 ( .A(n368), .Z(n1578) );
  IVSVTX4 U1629 ( .A(n1175), .Z(n1181) );
  AO6SVTX4 U1630 ( .A(n446), .B(n1574), .C(n1573), .Z(n1575) );
  ND2SVTX4 U1631 ( .A(n1201), .B(n824), .Z(n1266) );
  AO7ABSVTX8 U1632 ( .A(n1365), .B(n846), .C(n1474), .Z(n1506) );
  NR2ASVTX6 U1633 ( .A(n1232), .B(n1347), .Z(n1410) );
  IVSVTX4 U1634 ( .A(n1059), .Z(n1060) );
  IVSVTX10 U1635 ( .A(n813), .Z(n1688) );
  AO7SVTX8 U1636 ( .A(n1693), .B(n1689), .C(n1690), .Z(n1643) );
  IVSVTX4 U1637 ( .A(n919), .Z(n892) );
  IVSVTX2 U1638 ( .A(n1192), .Z(n1193) );
  IVSVTX2 U1639 ( .A(n1296), .Z(n1299) );
  ND2SVTX2 U1640 ( .A(n1626), .B(n1244), .Z(n1240) );
  IVSVTX4 U1641 ( .A(n874), .Z(n846) );
  IVSVTX2 U1642 ( .A(n1637), .Z(n1628) );
  ND3SVTX4 U1643 ( .A(n1431), .B(n873), .C(n1430), .Z(n1459) );
  IVSVTX2 U1644 ( .A(n1385), .Z(n1386) );
  IVSVTX2 U1645 ( .A(n383), .Z(n973) );
  NR2SVTX2 U1646 ( .A(n1270), .B(n1248), .Z(n1272) );
  IVSVTX2 U1647 ( .A(n1269), .Z(n1273) );
  IVSVTX4 U1648 ( .A(n1176), .Z(n1180) );
  IVSVTX2 U1649 ( .A(n297), .Z(n831) );
  ND3ABSVTX2 U1650 ( .A(N[4]), .B(N[5]), .C(N[2]), .Z(n926) );
  NR3SVTX2 U1651 ( .A(N[20]), .B(N[22]), .C(N[21]), .Z(n894) );
  F_ND2ASVTX2 U1652 ( .A(n1312), .B(n840), .Z(n1313) );
  ND2SVTX4 U1653 ( .A(n858), .B(n660), .Z(n1469) );
  NR2SVTX2 U1654 ( .A(n1823), .B(n1297), .Z(n1298) );
  IVSVTX2 U1655 ( .A(n1135), .Z(n1139) );
  ND2SVTX2 U1656 ( .A(n841), .B(n1163), .Z(n940) );
  F_AN2SVTX2 U1657 ( .A(n1625), .B(n1601), .Z(n1581) );
  ND2SVTX2 U1658 ( .A(n1232), .B(n282), .Z(n1372) );
  B_ND2SVTX1 U1659 ( .A(n1802), .B(n1801), .Z(n1807) );
  F_ND2SVTX1 U1660 ( .A(n1763), .B(n526), .Z(n1766) );
  ND2SVTX4 U1661 ( .A(n1382), .B(n1381), .Z(n1406) );
  ND2SVTX2 U1662 ( .A(O[27]), .B(n1332), .Z(n1333) );
  IVSVTX12 U1663 ( .A(n1232), .Z(n1823) );
  NR2ASVTX2 U1664 ( .A(n258), .B(n474), .Z(n1559) );
  ND2SVTX2 U1665 ( .A(n1625), .B(n474), .Z(n1548) );
  ND3ABSVTX6 U1666 ( .A(n1365), .B(n1317), .C(n1334), .Z(n1348) );
  NR2ASVTX2 U1667 ( .A(n1205), .B(n1118), .Z(n1171) );
  ND3ABSVTX2 U1668 ( .A(n1406), .B(n837), .C(n1394), .Z(n1385) );
  ND3SVTX1 U1669 ( .A(n544), .B(n1365), .C(N[3]), .Z(n1431) );
  AO7SVTX8 U1670 ( .A(n1531), .B(n1737), .C(n1734), .Z(n822) );
  EOSVTX4 U1671 ( .A(n1741), .B(n1740), .Z(O[13]) );
  ND2SVTX4 U1672 ( .A(n1020), .B(n1163), .Z(n1149) );
  ND2SVTX2 U1673 ( .A(n1134), .B(n1163), .Z(n1135) );
  AO2NSVTX4 U1674 ( .A(n1369), .B(O[27]), .C(n1368), .D(n232), .Z(n871) );
  AO2SVTX4 U1675 ( .A(n654), .B(n1176), .C(n1175), .D(n292), .Z(n824) );
  F_ND2SVTX1 U1676 ( .A(n1749), .B(n1748), .Z(n1751) );
  ND2ASVTX8 U1677 ( .A(n1524), .B(n1511), .Z(n1735) );
  NR3ASVTX2 U1678 ( .A(n959), .B(n1007), .C(n1150), .Z(n1153) );
  MUX21NSVTX2 U1679 ( .A(n827), .B(n1393), .S(n391), .Z(n1416) );
  ND2ASVTX8 U1680 ( .A(n483), .B(n1505), .Z(n1528) );
  IVSVTX2 U1681 ( .A(n1306), .Z(n1309) );
  AO7ABSVTX8 U1682 ( .A(n1062), .B(n728), .C(n1061), .Z(n1090) );
  OR2BSVTX4 U1683 ( .A(n267), .B(n1243), .Z(n1625) );
  NR2ASVTX6 U1684 ( .A(n1493), .B(n1602), .Z(n1304) );
  IVSVTX4 U1685 ( .A(n901), .Z(n844) );
  NR2SVTX4 U1686 ( .A(n1471), .B(n1470), .Z(n1472) );
  OR2SVTX8 U1687 ( .A(n1365), .B(n1480), .Z(n876) );
  AO4ABSVTX4 U1688 ( .C(n1183), .D(n1206), .A(n412), .B(n1175), .Z(n1220) );
  ND3SVTX4 U1689 ( .A(n1152), .B(n1151), .C(n1153), .Z(n1154) );
  ND3SVTX8 U1690 ( .A(n1237), .B(n1665), .C(n1238), .Z(n1246) );
  EOSVTX4 U1691 ( .A(n1715), .B(n1714), .Z(O[11]) );
  ND2ASVTX8 U1692 ( .A(n283), .B(n1525), .Z(n1737) );
  CTBUFSVTX8 U1693 ( .A(n1823), .Z(n833) );
  AN2SVTX4 U1694 ( .A(N[21]), .B(n906), .Z(n834) );
  AN2SVTX4 U1695 ( .A(n1379), .B(n863), .Z(n1331) );
  ND2SVTX4 U1696 ( .A(n1103), .B(n917), .Z(n836) );
  NR2SVTX4 U1697 ( .A(N[23]), .B(N[22]), .Z(n887) );
  AO2SVTX2 U1698 ( .A(n1232), .B(n1459), .C(n820), .D(n264), .Z(n1449) );
  ND4ABSVTX4 U1699 ( .A(N[18]), .B(N[30]), .C(n1013), .D(n881), .Z(n912) );
  ND2SVTX4 U1700 ( .A(n1408), .B(n1407), .Z(n1756) );
  IVSVTX0H U1701 ( .A(n1689), .Z(n1691) );
  ND3SVTX8 U1702 ( .A(n1413), .B(n1361), .C(n1411), .Z(n1767) );
  AO7NSVTX4 U1703 ( .A(n917), .B(n739), .C(n929), .Z(n850) );
  NR2ASVTX4 U1704 ( .A(n941), .B(n1033), .Z(n1036) );
  NR3SVTX8 U1705 ( .A(n705), .B(n964), .C(n965), .Z(n976) );
  IVSVTX2 U1706 ( .A(n930), .Z(n851) );
  IVSVTX2 U1707 ( .A(N[30]), .Z(n930) );
  ND2SVTX2 U1708 ( .A(n997), .B(n686), .Z(n991) );
  NR3SVTX4 U1709 ( .A(n1475), .B(n1048), .C(n1321), .Z(n1325) );
  ND3ABSVTX4 U1710 ( .A(n1130), .B(n1287), .C(n1286), .Z(n1488) );
  ND2SVTX4 U1711 ( .A(n1253), .B(n1252), .Z(n1269) );
  AO7SVTX6 U1712 ( .A(n1481), .B(n862), .C(n876), .Z(n1489) );
  NR3SVTX6 U1713 ( .A(n1375), .B(n1077), .C(n1067), .Z(n1088) );
  OR2SVTX2 U1714 ( .A(n1479), .B(n1478), .Z(n862) );
  NR2SVTX2 U1715 ( .A(n297), .B(n1006), .Z(n989) );
  NR2SVTX2 U1716 ( .A(n1345), .B(n282), .Z(n1353) );
  IVSVTX4 U1717 ( .A(n1338), .Z(n1339) );
  ND2SVTX2 U1718 ( .A(n1120), .B(n1119), .Z(n1124) );
  AO6ASVTX4 U1719 ( .A(n1110), .B(n1119), .C(n1109), .Z(n1114) );
  ND2SVTX4 U1720 ( .A(n1020), .B(n1119), .Z(n1021) );
  ND2SVTX2 U1721 ( .A(n1184), .B(n952), .Z(n1111) );
  AO7ASVTX4 U1722 ( .A(n1144), .B(n1030), .C(n295), .Z(n1146) );
  IVSVTX4 U1723 ( .A(n1427), .Z(n1003) );
  NR2SVTX2 U1724 ( .A(n1244), .B(n483), .Z(n1209) );
  ND3SVTX8 U1725 ( .A(n925), .B(n934), .C(n1041), .Z(n915) );
  AO6CSVTX8 U1726 ( .A(n1688), .B(n810), .C(n1649), .Z(n1677) );
  IVSVTX4 U1727 ( .A(n1675), .Z(n1649) );
  ND2SVTX4 U1728 ( .A(n1753), .B(n1600), .Z(n1603) );
  AN2SVTX4 U1729 ( .A(n1551), .B(n1550), .Z(n870) );
  ND3SVTX2 U1730 ( .A(N[1]), .B(n860), .C(n1029), .Z(n956) );
  NR2SVTX2 U1731 ( .A(n1572), .B(n1570), .Z(n1574) );
  AO6CSVTX8 U1732 ( .A(n1688), .B(n1686), .C(n1683), .Z(n1684) );
  AO6CSVTX2 U1733 ( .A(n1163), .B(n1162), .C(n930), .Z(n1164) );
  NR3ABSVTX2 U1734 ( .A(n1665), .B(n591), .C(n747), .Z(n1215) );
  ND3ASVTX8 U1735 ( .A(n1529), .B(n1528), .C(n1527), .Z(n1530) );
  IVSVTX2 U1736 ( .A(n1558), .Z(n1565) );
  ND2ASVTX8 U1737 ( .A(n393), .B(n1517), .Z(n1749) );
  ND2SVTX4 U1738 ( .A(n654), .B(n470), .Z(n1318) );
  ND2SVTX2 U1739 ( .A(n1440), .B(n1441), .Z(n1457) );
  NR2SVTX2 U1740 ( .A(n1409), .B(n1410), .Z(n1361) );
  IVSVTX2 U1741 ( .A(n1410), .Z(n1412) );
  ND2SVTX2 U1742 ( .A(n953), .B(n1029), .Z(n955) );
  NR2SVTX2 U1743 ( .A(n1335), .B(n710), .Z(n1336) );
  OR2SVTX4 U1744 ( .A(n1374), .B(n1068), .Z(n864) );
  AO7NSVTX4 U1745 ( .A(n1107), .B(n1830), .C(n954), .Z(n866) );
  AN2SVTX4 U1746 ( .A(n1484), .B(n1307), .Z(n867) );
  IVSVTX2 U1747 ( .A(n1742), .Z(n1736) );
  OR2SVTX2 U1748 ( .A(n276), .B(n1604), .Z(n877) );
  IVSVTX4 U1749 ( .A(n889), .Z(n1160) );
  NR3SVTX8 U1750 ( .A(N[23]), .B(N[22]), .C(N[25]), .Z(n881) );
  NR2SVTX8 U1751 ( .A(n914), .B(n885), .Z(n888) );
  ND2SVTX6 U1752 ( .A(n887), .B(n1013), .Z(n928) );
  ND2SVTX4 U1753 ( .A(n962), .B(n605), .Z(n904) );
  ND2SVTX8 U1754 ( .A(n901), .B(n923), .Z(n925) );
  IVSVTX8 U1755 ( .A(n925), .Z(n910) );
  ND2ASVTX8 U1756 ( .A(n912), .B(n910), .Z(n902) );
  IVSVTX2 U1757 ( .A(N[22]), .Z(n906) );
  IVSVTX4 U1758 ( .A(N[10]), .Z(n1015) );
  NR2SVTX4 U1759 ( .A(n928), .B(n294), .Z(n933) );
  NR3ABSVTX8 U1760 ( .A(N[0]), .B(n860), .C(n825), .Z(n1136) );
  IVSVTX0H U1761 ( .A(n1025), .Z(n946) );
  BFSVTX1 U1762 ( .A(N[11]), .Z(n1101) );
  BFSVTX1 U1763 ( .A(N[23]), .Z(n1191) );
  BFSVTX1 U1764 ( .A(N[15]), .Z(n1020) );
  ND2SVTX4 U1765 ( .A(n1149), .B(n1148), .Z(n1205) );
  ND2ASVTX8 U1766 ( .A(n975), .B(n974), .Z(n1550) );
  ND2ASVTX8 U1767 ( .A(n528), .B(n987), .Z(n992) );
  NR3ABSVTX8 U1768 ( .A(N[4]), .B(n1830), .C(n1030), .Z(n1097) );
  IVSVTX0H U1769 ( .A(n1013), .Z(n1014) );
  ND2SVTX2 U1770 ( .A(N[2]), .B(n1014), .Z(n1016) );
  ND2SVTX4 U1771 ( .A(n841), .B(n1119), .Z(n1018) );
  ND3SVTX2 U1772 ( .A(n941), .B(n1184), .C(n1065), .Z(n1022) );
  ND2ASVTX4 U1773 ( .A(n232), .B(n1308), .Z(n1039) );
  NR2SVTX2 U1774 ( .A(n1097), .B(n1008), .Z(n1034) );
  ND2ASVTX8 U1775 ( .A(n297), .B(n1163), .Z(n1056) );
  ND3SVTX8 U1776 ( .A(n1053), .B(n1054), .C(n1052), .Z(n1500) );
  NR2SVTX8 U1777 ( .A(n1500), .B(n1499), .Z(n1513) );
  ND3ASVTX8 U1778 ( .A(n298), .B(n850), .C(n688), .Z(n1064) );
  NR2SVTX6 U1779 ( .A(n1085), .B(n392), .Z(n1086) );
  IVSVTX2 U1780 ( .A(n1097), .Z(n1098) );
  NR2ASVTX6 U1781 ( .A(n1105), .B(n1104), .Z(n1206) );
  IVSVTX4 U1782 ( .A(n1108), .Z(n1109) );
  ND2SVTX4 U1783 ( .A(n1115), .B(n1114), .Z(n1199) );
  IVSVTX2 U1784 ( .A(n1113), .Z(n1117) );
  ND2SVTX2 U1785 ( .A(n524), .B(n1163), .Z(n1123) );
  NR2SVTX4 U1786 ( .A(n270), .B(n1125), .Z(n1478) );
  IVSVTX4 U1787 ( .A(n1376), .Z(n1129) );
  NR2SVTX8 U1788 ( .A(n1133), .B(n1132), .Z(n1468) );
  NR2SVTX4 U1789 ( .A(n1214), .B(n450), .Z(n1236) );
  NR2ASVTX6 U1790 ( .A(n1172), .B(n1171), .Z(n1189) );
  IVSVTX2 U1791 ( .A(n1220), .Z(n1173) );
  NR2SVTX8 U1792 ( .A(n1251), .B(n1291), .Z(n1277) );
  NR2ASVTX2 U1793 ( .A(n1191), .B(n1450), .Z(n1192) );
  AO7ABSVTX4 U1794 ( .A(n412), .B(n269), .C(n1196), .Z(n1221) );
  ND2SVTX4 U1795 ( .A(n1203), .B(n1466), .Z(n1262) );
  BFSVTX1 U1796 ( .A(n1247), .Z(n1218) );
  MUX21NSVTX2 U1797 ( .A(n1251), .B(n1222), .S(O[27]), .Z(n1223) );
  F_AN2SVTX2 U1798 ( .A(n1244), .B(n379), .Z(n1234) );
  IVSVTX4 U1799 ( .A(n1238), .Z(n1239) );
  F_ENSVTX2 U1800 ( .A(n1242), .B(n1551), .Z(n1564) );
  ND2SVTX4 U1802 ( .A(n1466), .B(n1264), .Z(n1253) );
  ND2SVTX4 U1803 ( .A(n1475), .B(n1251), .Z(n1252) );
  ND2SVTX4 U1804 ( .A(O[27]), .B(n1264), .Z(n1265) );
  AO7ABSVTX4 U1805 ( .A(n1466), .B(n1266), .C(n1265), .Z(n1268) );
  NR2ASVTX6 U1806 ( .A(n285), .B(n1268), .Z(n1297) );
  IVSVTX4 U1807 ( .A(n1268), .Z(n1271) );
  ND2SVTX4 U1808 ( .A(n1604), .B(n1602), .Z(n1300) );
  NR2SVTX2 U1809 ( .A(n287), .B(n1351), .Z(n1343) );
  NR2SVTX4 U1810 ( .A(n290), .B(n1310), .Z(n1328) );
  ND2ASVTX8 U1811 ( .A(n1316), .B(n1315), .Z(n1345) );
  NR2SVTX8 U1812 ( .A(n1320), .B(n1319), .Z(n1334) );
  ND2SVTX4 U1813 ( .A(n1051), .B(n1339), .Z(n1323) );
  IVSVTX4 U1814 ( .A(n1323), .Z(n1324) );
  ND2SVTX6 U1815 ( .A(n1358), .B(n1359), .Z(n1373) );
  IVSVTX4 U1816 ( .A(n1373), .Z(n1360) );
  IVSVTX2 U1817 ( .A(n1380), .Z(n1381) );
  ND2SVTX6 U1818 ( .A(n1399), .B(n1400), .Z(n1395) );
  NR3ABSVTX8 U1819 ( .A(n262), .B(n740), .C(n1437), .Z(n1396) );
  ENSVTX8 U1820 ( .A(n1405), .B(n1396), .Z(n1439) );
  ND2SVTX2 U1821 ( .A(n1432), .B(n1433), .Z(n1462) );
  ND2SVTX4 U1822 ( .A(n246), .B(n248), .Z(n1446) );
  ND2SVTX4 U1823 ( .A(n1459), .B(n1458), .Z(n1804) );
  ND2SVTX4 U1824 ( .A(n580), .B(n1502), .Z(n1533) );
  IVSVTX2 U1825 ( .A(n1476), .Z(n1477) );
  ND2SVTX4 U1826 ( .A(n1506), .B(n1489), .Z(n1487) );
  ND4ABSVTX8 U1827 ( .A(n579), .B(n1500), .C(n1502), .D(n1485), .Z(n1486) );
  NR2SVTX6 U1828 ( .A(n1728), .B(n1721), .Z(n1537) );
  NR2SVTX4 U1829 ( .A(n1823), .B(n1495), .Z(n1529) );
  ND2SVTX8 U1830 ( .A(n1497), .B(n1498), .Z(n1514) );
  ND4ABSVTX8 U1831 ( .A(n1529), .B(n1526), .C(n1528), .D(n1527), .Z(n1733) );
  ND2SVTX8 U1832 ( .A(n855), .B(n1735), .Z(n1532) );
  IVSVTX4 U1833 ( .A(n1522), .Z(n1517) );
  ND2SVTX6 U1834 ( .A(n1749), .B(n1710), .Z(n1743) );
  ND2ASVTX8 U1835 ( .A(n1518), .B(n1530), .Z(n1734) );
  AO17SVTX8 U1836 ( .A(n1540), .B(n1711), .C(n1539), .D(n1538), .Z(n1598) );
  ND3SVTX8 U1837 ( .A(n1541), .B(n1620), .C(n1598), .Z(n1542) );
  ND2SVTX6 U1838 ( .A(n1543), .B(n1542), .Z(n1544) );
  ENSVTX8 U1839 ( .A(n1237), .B(n1544), .Z(n1627) );
  ND2SVTX2 U1840 ( .A(n1581), .B(n1627), .Z(n1549) );
  F_ENSVTX2 U1841 ( .A(n1244), .B(n870), .Z(n1552) );
  ND2SVTX4 U1842 ( .A(n1554), .B(n1553), .Z(n1655) );
  NR2SVTX4 U1843 ( .A(n1554), .B(n1553), .Z(n1656) );
  IVSVTX0H U1844 ( .A(n1656), .Z(n1555) );
  ND2SVTX2 U1845 ( .A(n1655), .B(n1555), .Z(n1654) );
  IVSVTX4 U1846 ( .A(n1566), .Z(n1561) );
  FAS1SVTX4 U1847 ( .A(n1564), .B(1'b0), .CI(n1562), .CO(n1554), .Z(n1648) );
  EO3SVTX8 U1848 ( .A(n1558), .B(n861), .C(n1566), .Z(n1647) );
  HA1SVTX1 U1849 ( .A(n256), .B(n1567), .CO(n1556), .S(n1584) );
  BFSVTX2 U1850 ( .A(n1569), .Z(n1580) );
  NR2SVTX8 U1851 ( .A(n1646), .B(n1647), .Z(n1679) );
  AO7SVTX4 U1852 ( .A(n1572), .B(n685), .C(n1619), .Z(n1573) );
  AO7ABSVTX4 U1853 ( .A(n1632), .B(n1633), .C(n1582), .Z(n1645) );
  F_ENSVTX2 U1854 ( .A(n1584), .B(n1583), .Z(n1586) );
  IVSVTX2 U1855 ( .A(n1676), .Z(n1587) );
  ND2SVTX2 U1856 ( .A(n1589), .B(n1258), .Z(n1594) );
  ND2SVTX2 U1857 ( .A(n1257), .B(n1620), .Z(n1592) );
  F_ENSVTX2 U1858 ( .A(n1594), .B(n1593), .Z(n1595) );
  AN2BSVTX4 U1859 ( .A(n1595), .B(n1624), .Z(n1614) );
  ND2SVTX1 U1860 ( .A(n1599), .B(n1598), .Z(n1600) );
  FAS1SVTX4 U1861 ( .A(n1604), .B(n1603), .CI(n430), .CO(n1634), .Z(n1612) );
  NR2SVTX4 U1862 ( .A(n1612), .B(n1611), .Z(n1704) );
  F_ND2SVTX0H U1863 ( .A(n1257), .B(n229), .Z(n1609) );
  ND2SVTX4 U1864 ( .A(n1612), .B(n1611), .Z(n1705) );
  ND2SVTX4 U1865 ( .A(n275), .B(n1628), .Z(n1629) );
  NR2SVTX8 U1866 ( .A(n1642), .B(n1641), .Z(n1689) );
  NR2SVTX8 U1867 ( .A(n1639), .B(n1640), .Z(n1696) );
  NR2SVTX6 U1868 ( .A(n1689), .B(n1696), .Z(n1644) );
  AO6SVTX8 U1869 ( .A(n1688), .B(n1652), .C(n1651), .Z(n1653) );
  EOSVTX8 U1870 ( .A(n1654), .B(n1653), .Z(O[24]) );
  NR2SVTX4 U1871 ( .A(n1672), .B(n1656), .Z(n1658) );
  ND2SVTX4 U1872 ( .A(n1658), .B(n1676), .Z(n1661) );
  IVSVTX2 U1873 ( .A(n1824), .Z(n1671) );
  IVSVTX0H U1874 ( .A(n1672), .Z(n1673) );
  ND2SVTX2 U1875 ( .A(n1674), .B(n1673), .Z(n1678) );
  EOSVTX8 U1876 ( .A(n1678), .B(n1677), .Z(O[23]) );
  IVSVTX0H U1877 ( .A(n1679), .Z(n1681) );
  ND2SVTX2 U1878 ( .A(n1681), .B(n1680), .Z(n1685) );
  EOSVTX8 U1879 ( .A(n1685), .B(n1684), .Z(O[22]) );
  ND2SVTX2 U1880 ( .A(n1686), .B(n1683), .Z(n1687) );
  ND2SVTX2 U1881 ( .A(n1691), .B(n1690), .Z(n1695) );
  ND2SVTX4 U1882 ( .A(n854), .B(n1697), .Z(n1698) );
  ND2SVTX2 U1883 ( .A(n1706), .B(n1705), .Z(n1707) );
  ENSVTX4 U1884 ( .A(n1708), .B(n1707), .Z(O[17]) );
  IVSVTX2 U1885 ( .A(n1711), .Z(n1712) );
  BFSVTX1 U1886 ( .A(n1718), .Z(n1726) );
  IVSVTX0H U1887 ( .A(n1726), .Z(n1727) );
  AO7SVTX1 U1888 ( .A(n370), .B(n1727), .C(n1716), .Z(n1729) );
  NR2SVTX2 U1889 ( .A(n1736), .B(n1743), .Z(n1739) );
  AO7SVTX1 U1890 ( .A(n495), .B(n1736), .C(n396), .Z(n1738) );
  BFSVTX4 U1891 ( .A(n1755), .Z(n1772) );
  BFSVTX4 U1892 ( .A(n1757), .Z(n1758) );
  AO7SVTX2 U1893 ( .A(n1793), .B(n238), .C(n431), .Z(n1760) );
  AO7SVTX2 U1894 ( .A(n1793), .B(n1792), .C(n1764), .Z(n1765) );
  F_ND2SVTX1 U1895 ( .A(n1768), .B(n1767), .Z(n1777) );
  IVSVTX1 U1896 ( .A(n238), .Z(n1769) );
  AO6SVTX1 U1897 ( .A(n1773), .B(n1772), .C(n1771), .Z(n1774) );
  AO7SVTX2 U1898 ( .A(n1793), .B(n1775), .C(n1774), .Z(n1776) );
  ND2SVTX2 U1899 ( .A(n1779), .B(n1780), .Z(n1786) );
  AO6SVTX1 U1900 ( .A(n406), .B(n346), .C(n1782), .Z(n1783) );
  AO7SVTX2 U1901 ( .A(n1784), .B(n1793), .C(n1783), .Z(n1785) );
  AO7SVTX2 U1902 ( .A(n1418), .B(n1793), .C(n1789), .Z(n1790) );
  BFSVTX4 U1903 ( .A(n1795), .Z(n1816) );
  AO6SVTX1 U1904 ( .A(n429), .B(n1811), .C(n312), .Z(n1798) );
  IVSVTX2 U1905 ( .A(n1803), .Z(n1821) );
  NR2SVTX2 U1906 ( .A(n1816), .B(n1812), .Z(n1818) );
  AO7SVTX1 U1907 ( .A(n1816), .B(n1815), .C(n1814), .Z(n1817) );
  AO7SVTX1 U1908 ( .A(n819), .B(n258), .C(n1823), .Z(n1825) );
  ND2SVTX2 U1909 ( .A(n1825), .B(n1824), .Z(n1826) );
  EOSVTX8 U1910 ( .A(n1829), .B(n1828), .Z(O[26]) );
endmodule

