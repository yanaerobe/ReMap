
module remap ( m1, m2 );
  input [27:0] m1;
  output [26:0] m2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787;

  IVSVTX0H U3 ( .A(n657), .Z(n754) );
  IVSVTX0H U4 ( .A(n699), .Z(n761) );
  IVSVTX0H U5 ( .A(n650), .Z(n665) );
  AO6SVTX6 U6 ( .A(n786), .B(n784), .C(n740), .Z(n747) );
  AO11NSVTX1 U7 ( .A(n388), .B(n720), .C(n719), .D(n718), .E(n717), .F(m1[21]), 
        .Z(n735) );
  AO11NSVTX1 U8 ( .A(n388), .B(n238), .C(n719), .D(n237), .E(n717), .F(m1[20]), 
        .Z(n714) );
  IVSVTX0H U9 ( .A(n776), .Z(n717) );
  FA1SVTX1 U10 ( .A(m1[21]), .B(n321), .CI(n320), .CO(n240), .Z(n591) );
  FA1SVTX1 U11 ( .A(m1[13]), .B(n437), .CI(n546), .CO(n571), .Z(n566) );
  FA1SVTX1 U12 ( .A(m1[4]), .B(n470), .CI(n546), .CO(n521), .Z(n518) );
  F_FA1SVTX1 U13 ( .A(m1[7]), .B(n544), .CI(n546), .CO(n553), .Z(n550) );
  F_FA1SVTX1 U14 ( .A(m1[8]), .B(n533), .CI(n546), .CO(n555), .Z(n552) );
  F_FA1SVTX1 U15 ( .A(m1[15]), .B(n427), .CI(n546), .CO(n575), .Z(n572) );
  F_FA1SVTX1 U16 ( .A(n401), .B(n387), .CI(n386), .CO(n587), .Z(n584) );
  FA1SVTX4 U17 ( .A(m1[19]), .B(n376), .CI(n375), .CO(n590), .Z(n586) );
  FA1SVTX2 U18 ( .A(n324), .B(n399), .CI(n398), .CO(n585), .Z(n576) );
  F_FA1SVTX1 U19 ( .A(m1[5]), .B(n545), .CI(n546), .CO(n549), .Z(n520) );
  ND4SVTX1 U20 ( .A(n420), .B(n397), .C(n485), .D(n396), .Z(n421) );
  AO11NSVTX1 U21 ( .A(n543), .B(n392), .C(n719), .D(n391), .E(n540), .F(m1[14]), .Z(n422) );
  IVSVTX0H U22 ( .A(n713), .Z(n727) );
  AO6NSVTX1 U23 ( .A(n505), .B(n504), .C(n503), .Z(n771) );
  ND4SVTX1 U24 ( .A(n482), .B(n481), .C(n495), .D(n480), .Z(n512) );
  NR4ABCSVTX1 U25 ( .A(n497), .B(n373), .C(n397), .D(n721), .Z(n480) );
  IVSVTX0H U26 ( .A(n405), .Z(n418) );
  NR2ASVTX1 U27 ( .A(n373), .B(n367), .Z(n260) );
  F_MUX21NSVTX0H U28 ( .A(n357), .B(m1[24]), .S(n262), .Z(n147) );
  NR2ASVTX1 U29 ( .A(n293), .B(n315), .Z(n301) );
  ND4SVTX1 U30 ( .A(n352), .B(n314), .C(n329), .D(n353), .Z(n205) );
  IVSVTX0H U31 ( .A(n357), .Z(n283) );
  IVSVTX0H U32 ( .A(n73), .Z(n258) );
  NR2ASVTX1 U33 ( .A(n295), .B(n120), .Z(n248) );
  AO7SVTX1 U34 ( .A(n90), .B(n215), .C(n123), .Z(n114) );
  IVSVTX0H U35 ( .A(n273), .Z(n266) );
  IVSVTX0H U36 ( .A(m1[27]), .Z(n108) );
  IVSVTX2 U37 ( .A(n311), .Z(n297) );
  IVSVTX0H U38 ( .A(n327), .Z(n293) );
  IVSVTX0H U39 ( .A(n123), .Z(n119) );
  IVSVTX0H U40 ( .A(n124), .Z(n90) );
  AO21SVTX1 U41 ( .A(n163), .B(n8), .C(n7), .D(m1[11]), .Z(n9) );
  IVSVTX2 U42 ( .A(m1[23]), .Z(n295) );
  IVSVTX2 U43 ( .A(m1[10]), .Z(n134) );
  B_ND2SVTX0H U44 ( .A(n197), .B(n196), .Z(n198) );
  ND2ASVTX1 U45 ( .A(n39), .B(m1[2]), .Z(n40) );
  IVSVTX0H U46 ( .A(n180), .Z(n181) );
  B_ND2SVTX0H U47 ( .A(m1[8]), .B(m1[9]), .Z(n194) );
  ND2ASVTX1 U48 ( .A(m1[23]), .B(n706), .Z(n256) );
  B_ND2SVTX0H U49 ( .A(m1[20]), .B(n252), .Z(n270) );
  B_ND2SVTX0H U50 ( .A(n311), .B(n271), .Z(n224) );
  ND2ASVTX1 U51 ( .A(m1[11]), .B(n81), .Z(n187) );
  AO17SVTX1 U52 ( .A(n81), .B(n75), .C(n167), .D(n184), .Z(n56) );
  AO1ABSVTX2 U53 ( .A(n324), .B(m1[19]), .C(n354), .D(n149), .Z(n116) );
  F_ND2SVTX0H U54 ( .A(n476), .B(n456), .Z(n453) );
  F_ND2SVTX0H U55 ( .A(n481), .B(n291), .Z(n393) );
  NR3SVTX1 U56 ( .A(n285), .B(n284), .C(n283), .Z(n363) );
  NR3SVTX1 U57 ( .A(n395), .B(n394), .C(n393), .Z(n420) );
  NR4SVTX1 U58 ( .A(n344), .B(n366), .C(n343), .D(n342), .Z(n396) );
  ND2ASVTX1 U59 ( .A(n273), .B(n147), .Z(n316) );
  IVSVTX0H U60 ( .A(n614), .Z(n618) );
  AO7SVTX6 U61 ( .A(n749), .B(n752), .C(n751), .Z(n786) );
  ENSVTX0H U62 ( .A(n596), .B(n731), .Z(m2[21]) );
  EOSVTX0H U63 ( .A(n604), .B(n681), .Z(m2[7]) );
  AO6SVTX6 U64 ( .A(n583), .B(n598), .C(n582), .Z(n624) );
  AO6SVTX4 U65 ( .A(n523), .B(n699), .C(n522), .Z(n601) );
  CTIVSVTX2 U66 ( .A(n662), .Z(n640) );
  B_ND2SVTX1 U67 ( .A(n671), .B(n670), .Z(n676) );
  F_IVSVTX1 U68 ( .A(n769), .Z(n508) );
  B_ND2SVTX1 U69 ( .A(n779), .B(n778), .Z(n783) );
  AO11NSVTX2 U70 ( .A(n543), .B(n351), .C(n719), .D(n350), .E(n540), .F(m1[16]), .Z(n387) );
  ND3SVTX2 U71 ( .A(n501), .B(n374), .C(n480), .Z(n386) );
  AO7SVTX2 U72 ( .A(n362), .B(n361), .C(n360), .Z(n394) );
  F_IVSVTX1 U73 ( .A(n34), .Z(n30) );
  B_ND2SVTX2 U74 ( .A(n334), .B(n333), .Z(n407) );
  ND4SVTX2 U75 ( .A(m1[26]), .B(m1[20]), .C(n324), .D(n19), .Z(n34) );
  F_IVSVTX1 U76 ( .A(n64), .Z(n12) );
  IVSVTX2 U77 ( .A(n272), .Z(n296) );
  AO17SVTX2 U78 ( .A(m1[9]), .B(n26), .C(n25), .D(n24), .Z(n28) );
  B_ND2SVTX2 U79 ( .A(m1[23]), .B(n120), .Z(n213) );
  CTIVSVTX4 U80 ( .A(m1[20]), .Z(n149) );
  IVSVTX2 U81 ( .A(n785), .Z(n740) );
  EOSVTX0H U82 ( .A(n767), .B(n766), .Z(m2[2]) );
  AO7SVTX4 U83 ( .A(n767), .B(n763), .C(n765), .Z(n699) );
  FA1SVTX2 U84 ( .A(m1[22]), .B(n714), .CI(n713), .CO(n733), .Z(n239) );
  B_ND2SVTX2 U85 ( .A(n639), .B(n638), .Z(n642) );
  AO6SVTX4 U86 ( .A(n702), .B(n705), .C(n511), .Z(n767) );
  B_ND2SVTX1 U87 ( .A(n666), .B(n665), .Z(n668) );
  B_ND2SVTX1 U88 ( .A(n672), .B(n597), .Z(n599) );
  EOSVTX0H U89 ( .A(m1[24]), .B(n716), .Z(n237) );
  B_ND2SVTX1 U90 ( .A(n607), .B(n606), .Z(n617) );
  B_ND2SVTX2 U91 ( .A(n295), .B(n236), .Z(n716) );
  B_ND2SVTX2 U92 ( .A(n742), .B(n741), .Z(n746) );
  BFSVTX6 U93 ( .A(n388), .Z(n543) );
  B_ND2SVTX2 U94 ( .A(n487), .B(n727), .Z(n736) );
  NR3ABSVTX4 U95 ( .A(n345), .B(n289), .C(n69), .Z(n487) );
  NR2ASVTX2 U96 ( .A(n726), .B(n344), .Z(n317) );
  ND4ABCSVTX2 U97 ( .A(n290), .B(n339), .C(n367), .D(n382), .Z(n479) );
  AO1ABSVTX1 U98 ( .A(n287), .B(n333), .C(n286), .D(n363), .Z(n288) );
  B_ND2SVTX0H U99 ( .A(n293), .B(n297), .Z(n276) );
  AO21SVTX2 U100 ( .A(n275), .B(n296), .C(n274), .D(n273), .Z(n292) );
  CTIVSVTX2 U101 ( .A(n285), .Z(n106) );
  IVSVTX2 U102 ( .A(n265), .Z(n271) );
  B_ND2SVTX2 U103 ( .A(n324), .B(n191), .Z(n180) );
  B_ND2SVTX1 U104 ( .A(n169), .B(n167), .Z(n172) );
  IVSVTX2 U105 ( .A(n225), .Z(n268) );
  IVSVTX4 U106 ( .A(n72), .Z(n401) );
  IVSVTX2 U107 ( .A(m1[24]), .Z(n706) );
  IVSVTX4 U108 ( .A(m1[21]), .Z(n314) );
  AO6SVTX6 U109 ( .A(n731), .B(n730), .C(n729), .Z(n752) );
  IVSVTX4 U110 ( .A(n598), .Z(n673) );
  B_ND2SVTX1 U111 ( .A(n751), .B(n750), .Z(n753) );
  AO7SVTX6 U112 ( .A(n601), .B(n559), .C(n558), .Z(n598) );
  CTIVSVTX2 U113 ( .A(n728), .Z(n729) );
  B_ND2SVTX2 U114 ( .A(n728), .B(n730), .Z(n596) );
  NR2SVTX2 U115 ( .A(n733), .B(n732), .Z(n749) );
  B_ND2SVTX2 U116 ( .A(n739), .B(n738), .Z(n785) );
  B_ND2SVTX2 U117 ( .A(n623), .B(n622), .Z(n628) );
  B_ND2SVTX2 U118 ( .A(n638), .B(n1), .Z(n632) );
  B_ND2SVTX2 U119 ( .A(n587), .B(n586), .Z(n639) );
  B_ND2SVTX2 U120 ( .A(n619), .B(n618), .Z(n621) );
  AO6SVTX2 U121 ( .A(n569), .B(n647), .C(n568), .Z(n609) );
  NR2SVTX1 U122 ( .A(m1[24]), .B(n716), .Z(n718) );
  B_ND2SVTX2 U123 ( .A(n510), .B(n509), .Z(n703) );
  B_ND2SVTX2 U124 ( .A(n706), .B(n235), .Z(n715) );
  NR2SVTX1 U125 ( .A(n708), .B(n388), .Z(n774) );
  IVSVTX6 U126 ( .A(n489), .Z(n719) );
  B_ND2SVTX1 U127 ( .A(n410), .B(n412), .Z(n366) );
  F_AN2SVTX2 U128 ( .A(n108), .B(n126), .Z(n711) );
  B_ND2SVTX1 U129 ( .A(n332), .B(n331), .Z(n484) );
  NR4SVTX2 U130 ( .A(m1[23]), .B(n296), .C(n283), .D(n279), .Z(n333) );
  ND3SVTX2 U131 ( .A(n63), .B(n115), .C(n13), .Z(n14) );
  AO3SVTX2 U132 ( .A(n204), .B(n287), .C(n221), .D(n357), .Z(n280) );
  B_ND2SVTX1 U133 ( .A(m1[20]), .B(n297), .Z(n309) );
  CTIVSVTX2 U134 ( .A(n231), .Z(n281) );
  B_IVSVTX1 U135 ( .A(n15), .Z(n16) );
  B_ND2SVTX2 U136 ( .A(n106), .B(n105), .Z(n249) );
  NR3SVTX2 U137 ( .A(n59), .B(n47), .C(n153), .Z(n57) );
  CTIVSVTX2 U138 ( .A(n256), .Z(n105) );
  B_ND2SVTX1 U139 ( .A(n456), .B(n472), .Z(n467) );
  F_ND2ASVTX2 U140 ( .A(n295), .B(m1[20]), .Z(n231) );
  F_ND2ASVTX2 U141 ( .A(m1[22]), .B(n356), .Z(n120) );
  NR2ASVTX4 U142 ( .A(n706), .B(n273), .Z(n357) );
  B_ND2SVTX2 U143 ( .A(n184), .B(n75), .Z(n191) );
  B_ND2SVTX1 U144 ( .A(m1[19]), .B(n401), .Z(n143) );
  F_ND2SVTX1 U145 ( .A(n475), .B(n476), .Z(n455) );
  B_IVSVTX1 U146 ( .A(n40), .Z(n175) );
  AN2ABSVTX2 U147 ( .A(m1[26]), .B(m1[27]), .Z(n352) );
  F_ND2ASVTX2 U148 ( .A(m1[27]), .B(n115), .Z(n123) );
  IVSVTX2 U149 ( .A(m1[18]), .Z(n72) );
  B_ND2SVTX2 U150 ( .A(n78), .B(n179), .Z(n142) );
  CTIVSVTX2 U151 ( .A(m1[7]), .Z(n160) );
  EOSVTX0H U152 ( .A(n691), .B(n690), .Z(m2[6]) );
  EOSVTX0H U153 ( .A(n599), .B(n673), .Z(m2[9]) );
  AO7SVTX6 U154 ( .A(n595), .B(n624), .C(n594), .Z(n731) );
  B_ND2SVTX1 U155 ( .A(n785), .B(n784), .Z(n787) );
  EOSVTX0H U156 ( .A(n762), .B(n761), .Z(m2[3]) );
  B_ND2SVTX2 U157 ( .A(n240), .B(n239), .Z(n728) );
  B_ND2SVTX2 U158 ( .A(n733), .B(n732), .Z(n751) );
  F_ND2SVTX1 U159 ( .A(n631), .B(n630), .Z(n637) );
  OR2SVTX2 U160 ( .A(n592), .B(n591), .Z(n622) );
  B_ND2SVTX2 U161 ( .A(n592), .B(n591), .Z(n623) );
  F_ND2SVTX1 U162 ( .A(n765), .B(n764), .Z(n766) );
  B_ND2SVTX1 U163 ( .A(n656), .B(n655), .Z(n661) );
  B_ND2SVTX1 U164 ( .A(n703), .B(n702), .Z(n704) );
  B_ND2SVTX1 U165 ( .A(n645), .B(n644), .Z(n653) );
  B_ND2SVTX1 U166 ( .A(n698), .B(n697), .Z(n701) );
  B_ND2SVTX1 U167 ( .A(n760), .B(n759), .Z(n762) );
  IVSVTX2 U168 ( .A(n703), .Z(n511) );
  ND2SVTX2 U169 ( .A(n569), .B(n646), .Z(n610) );
  B_ND2SVTX1 U170 ( .A(n755), .B(n754), .Z(n757) );
  AO6SVTX2 U171 ( .A(n557), .B(n602), .C(n556), .Z(n558) );
  B_ND2SVTX1 U172 ( .A(n680), .B(n600), .Z(n604) );
  B_ND2SVTX1 U173 ( .A(n679), .B(n678), .Z(n684) );
  B_ND2SVTX2 U174 ( .A(n557), .B(n603), .Z(n559) );
  ND2SVTX2 U175 ( .A(n579), .B(n608), .Z(n581) );
  B_ND2SVTX1 U176 ( .A(n687), .B(n686), .Z(n691) );
  F_ND2SVTX1 U177 ( .A(n693), .B(n692), .Z(n695) );
  B_ND2SVTX1 U178 ( .A(n662), .B(n1), .Z(n664) );
  AO7SVTX2 U179 ( .A(n755), .B(n654), .C(n656), .Z(n611) );
  B_ND2SVTX1 U180 ( .A(n769), .B(n768), .Z(n770) );
  B_ND2SVTX2 U181 ( .A(n517), .B(n516), .Z(n765) );
  B_ND2SVTX1 U182 ( .A(n746), .B(n745), .Z(n748) );
  AO7SVTX2 U183 ( .A(n693), .B(n685), .C(n687), .Z(n602) );
  B_ND2SVTX2 U184 ( .A(n585), .B(n584), .Z(n662) );
  AO7SVTX2 U185 ( .A(n680), .B(n677), .C(n679), .Z(n556) );
  AO7SVTX2 U186 ( .A(n672), .B(n669), .C(n671), .Z(n647) );
  OR2SVTX2 U187 ( .A(n585), .B(n584), .Z(n1) );
  ND2SVTX2 U188 ( .A(n571), .B(n570), .Z(n755) );
  B_ND2SVTX2 U189 ( .A(n551), .B(n550), .Z(n687) );
  OR2SVTX2 U190 ( .A(n710), .B(n709), .Z(n781) );
  B_ND2SVTX2 U191 ( .A(n573), .B(n572), .Z(n656) );
  B_ND2SVTX2 U192 ( .A(n567), .B(n566), .Z(n645) );
  B_ND2SVTX2 U193 ( .A(n561), .B(n560), .Z(n672) );
  B_ND2SVTX2 U194 ( .A(n521), .B(n520), .Z(n698) );
  ND2SVTX2 U195 ( .A(n565), .B(n564), .Z(n666) );
  B_ND2SVTX2 U196 ( .A(n575), .B(n574), .Z(n619) );
  B_ND2SVTX2 U197 ( .A(n553), .B(n552), .Z(n680) );
  B_ND2SVTX2 U198 ( .A(n507), .B(n506), .Z(n769) );
  B_ND2SVTX2 U199 ( .A(n577), .B(n576), .Z(n607) );
  B_ND2SVTX2 U200 ( .A(n555), .B(n554), .Z(n679) );
  B_ND2SVTX2 U201 ( .A(n519), .B(n518), .Z(n760) );
  FAS1SVTX2 U202 ( .A(m1[16]), .B(n422), .CI(n421), .CO(n577), .Z(n574) );
  ND2SVTX2 U203 ( .A(n330), .B(n322), .Z(n241) );
  OR2SVTX2 U204 ( .A(n385), .B(n384), .Z(n398) );
  ND2SVTX2 U205 ( .A(n149), .B(n377), .Z(n348) );
  OR3SVTX2 U206 ( .A(n371), .B(n723), .C(n736), .Z(n320) );
  IVSVTX4 U207 ( .A(n776), .Z(n540) );
  NR4SVTX4 U208 ( .A(n418), .B(n417), .C(n490), .D(n416), .Z(n483) );
  NR3ABSVTX4 U209 ( .A(n283), .B(n316), .C(n479), .Z(n776) );
  B_ND2SVTX2 U210 ( .A(n72), .B(n400), .Z(n389) );
  AO17SVTX2 U211 ( .A(n255), .B(n31), .C(n30), .D(n29), .Z(n289) );
  ND4SVTX6 U212 ( .A(n405), .B(n383), .C(n497), .D(n127), .Z(n708) );
  ND3SVTX1 U213 ( .A(n341), .B(n415), .C(n340), .Z(n342) );
  NR2ASVTX4 U214 ( .A(n341), .B(n369), .Z(n383) );
  B_ND2SVTX2 U215 ( .A(n170), .B(n428), .Z(n423) );
  F_ND2SVTX1 U216 ( .A(n313), .B(n253), .Z(n372) );
  IVSVTX2 U217 ( .A(n711), .Z(n127) );
  AO1ABSVTX4 U218 ( .A(n273), .B(n262), .C(n357), .D(n158), .Z(n367) );
  AO6SVTX2 U219 ( .A(n218), .B(n245), .C(n266), .Z(n158) );
  F_IVSVTX1 U220 ( .A(n66), .Z(n29) );
  AO17SVTX1 U221 ( .A(n271), .B(n315), .C(n272), .D(n295), .Z(n220) );
  ND2SVTX2 U222 ( .A(n75), .B(n438), .Z(n433) );
  IVSVTX1 U223 ( .A(n362), .Z(n156) );
  IVSVTX2 U224 ( .A(n282), .Z(n155) );
  CTIVSVTX2 U225 ( .A(n17), .Z(n18) );
  F_ND2SVTX1 U226 ( .A(n111), .B(n110), .Z(n113) );
  AO3SVTX2 U227 ( .A(n58), .B(n68), .C(n57), .D(n60), .Z(n481) );
  B_ND2SVTX2 U228 ( .A(m1[21]), .B(n121), .Z(n89) );
  AO6SVTX2 U229 ( .A(n88), .B(n87), .C(n168), .Z(n121) );
  ND2SVTX2 U230 ( .A(n71), .B(n448), .Z(n443) );
  AO3SVTX2 U231 ( .A(n149), .B(n16), .C(n106), .D(n295), .Z(n31) );
  F_ND2SVTX1 U232 ( .A(n314), .B(n329), .Z(n189) );
  NR3SVTX6 U233 ( .A(n21), .B(n5), .C(n4), .Z(n311) );
  B_ND2SVTX2 U234 ( .A(n101), .B(n100), .Z(n111) );
  B_ND2SVTX2 U235 ( .A(m1[20]), .B(n293), .Z(n272) );
  NR2SVTX1 U236 ( .A(n327), .B(n271), .Z(n275) );
  F_ND2SVTX1 U237 ( .A(n11), .B(n354), .Z(n15) );
  AO17SVTX1 U238 ( .A(n166), .B(n20), .C(n199), .D(n179), .Z(n26) );
  AO7SVTX1 U239 ( .A(n99), .B(n98), .C(n184), .Z(n101) );
  ND2SVTX2 U240 ( .A(n134), .B(n529), .Z(n524) );
  B_ND2SVTX2 U241 ( .A(m1[22]), .B(m1[21]), .Z(n327) );
  B_ND2SVTX1 U242 ( .A(m1[22]), .B(m1[20]), .Z(n46) );
  NR3ABSVTX1 U243 ( .A(m1[8]), .B(m1[10]), .C(n199), .Z(n93) );
  B_ND2SVTX1 U244 ( .A(m1[19]), .B(n38), .Z(n65) );
  B_ND2SVTX2 U245 ( .A(n199), .B(n139), .Z(n5) );
  IVSVTX4 U246 ( .A(m1[15]), .Z(n184) );
  ND3SVTX1 U247 ( .A(n81), .B(n134), .C(n75), .Z(n86) );
  CTIVSVTX2 U248 ( .A(m1[16]), .Z(n170) );
  ND2ASVTX4 U249 ( .A(m1[25]), .B(n352), .Z(n273) );
  B_ND2SVTX2 U250 ( .A(n160), .B(n179), .Z(n534) );
  B_ND2SVTX2 U251 ( .A(m1[26]), .B(m1[25]), .Z(n115) );
  F_IVSVTX0H U252 ( .A(n233), .Z(n226) );
  AO6SVTX2 U253 ( .A(n174), .B(m1[4]), .C(m1[7]), .Z(n178) );
  ND3SVTX2 U254 ( .A(m1[19]), .B(m1[14]), .C(m1[15]), .Z(n133) );
  AO6SVTX2 U255 ( .A(n136), .B(n134), .C(n133), .Z(n135) );
  AO3SVTX1 U256 ( .A(m1[13]), .B(n187), .C(n135), .D(n401), .Z(n146) );
  NR2SVTX2 U257 ( .A(m1[5]), .B(m1[4]), .Z(n139) );
  F_ND2ASVTX2 U258 ( .A(m1[22]), .B(n314), .Z(n285) );
  AO7SVTX4 U259 ( .A(n629), .B(n633), .C(n631), .Z(n625) );
  FA1SVTX1 U260 ( .A(m1[10]), .B(n452), .CI(n546), .CO(n563), .Z(n560) );
  ND2SVTX2 U261 ( .A(m1[9]), .B(m1[10]), .Z(n176) );
  NR2SVTX2 U262 ( .A(m1[24]), .B(m1[27]), .Z(n124) );
  NR2ASVTX2 U263 ( .A(n412), .B(n411), .Z(n413) );
  NR2ASVTX2 U264 ( .A(m1[25]), .B(n311), .Z(n252) );
  NR2SVTX2 U265 ( .A(n355), .B(n272), .Z(n204) );
  ND2SVTX2 U266 ( .A(n456), .B(n454), .Z(n128) );
  NR2SVTX2 U267 ( .A(n152), .B(n221), .Z(n290) );
  AO7SVTX2 U268 ( .A(n75), .B(n18), .C(n184), .Z(n19) );
  NR3SVTX2 U269 ( .A(n179), .B(n6), .C(n200), .Z(n7) );
  NR2SVTX2 U270 ( .A(n137), .B(n515), .Z(n6) );
  IVSVTX2 U271 ( .A(n371), .Z(n492) );
  F_EOSVTX2 U272 ( .A(n617), .B(n616), .Z(m2[16]) );
  AO6SVTX2 U273 ( .A(n620), .B(n618), .C(n615), .Z(n616) );
  F_ND2ASVTX2 U274 ( .A(n297), .B(n33), .Z(n304) );
  NR2SVTX2 U275 ( .A(n455), .B(n128), .Z(n462) );
  EOSVTX2 U276 ( .A(n748), .B(n747), .Z(m2[24]) );
  NR3SVTX2 U277 ( .A(n32), .B(n180), .C(n231), .Z(n10) );
  F_ENSVTX2 U278 ( .A(n743), .B(n780), .Z(m2[25]) );
  IVSVTX2 U279 ( .A(m1[5]), .Z(n465) );
  EOSVTX4 U280 ( .A(n783), .B(n782), .Z(m2[26]) );
  AO20SVTX2 U281 ( .A(n456), .B(n166), .C(n165), .D(n164), .Z(n173) );
  ND2SVTX2 U282 ( .A(n129), .B(n462), .Z(n525) );
  NR2SVTX2 U283 ( .A(m1[13]), .B(n443), .Z(n438) );
  ND2SVTX4 U284 ( .A(n168), .B(n378), .Z(n349) );
  NR2SVTX2 U285 ( .A(n401), .B(n390), .Z(n378) );
  ND2SVTX4 U286 ( .A(n132), .B(n402), .Z(n390) );
  NR2SVTX2 U287 ( .A(m1[10]), .B(n525), .Z(n449) );
  ENSVTX2 U288 ( .A(n787), .B(n786), .Z(m2[23]) );
  ND4SVTX2 U289 ( .A(n410), .B(n481), .C(n373), .D(n495), .Z(n69) );
  NR2SVTX0H U290 ( .A(n356), .B(n355), .Z(n359) );
  AO17ASVTX2 U291 ( .A(n297), .B(n114), .C(n119), .D(n14), .Z(n345) );
  AO7SVTX1 U292 ( .A(m1[24]), .B(n12), .C(m1[26]), .Z(n13) );
  NR2SVTX0H U293 ( .A(m1[25]), .B(n715), .Z(n720) );
  AO7ABSVTX1 U294 ( .A(m1[1]), .B(m1[0]), .C(n488), .Z(n76) );
  AN2SVTX0H U295 ( .A(m1[5]), .B(m1[6]), .Z(n174) );
  NR3SVTX1 U296 ( .A(n163), .B(m1[5]), .C(m1[6]), .Z(n165) );
  AO20SVTX1 U297 ( .A(n465), .B(n456), .C(n199), .D(n179), .Z(n8) );
  AO20SVTX1 U298 ( .A(n269), .B(n268), .C(n267), .D(n266), .Z(n305) );
  AO20SVTX1 U299 ( .A(m1[10]), .B(n43), .C(m1[11]), .D(n42), .Z(n44) );
  F_ND2SVTX0H U300 ( .A(n130), .B(n170), .Z(n42) );
  F_ND2SVTX0H U301 ( .A(n471), .B(n454), .Z(n460) );
  AN2SVTX0H U302 ( .A(m1[25]), .B(m1[24]), .Z(n157) );
  NR2ASVTX1 U303 ( .A(n722), .B(n721), .Z(n725) );
  AO7SVTX2 U304 ( .A(n760), .B(n696), .C(n698), .Z(n522) );
  AO7SVTX2 U305 ( .A(n666), .B(n643), .C(n645), .Z(n568) );
  AN2SVTX0H U306 ( .A(m1[0]), .B(n502), .Z(n503) );
  NR2SVTX2 U307 ( .A(n551), .B(n550), .Z(n685) );
  F_IVSVTX0H U308 ( .A(n623), .Z(n593) );
  NR2SVTX0H U309 ( .A(m1[11]), .B(m1[13]), .Z(n96) );
  IVSVTX0H U310 ( .A(m1[9]), .Z(n78) );
  AO6CSVTX1 U311 ( .A(n465), .B(n48), .C(m1[7]), .Z(n77) );
  F_ND2SVTX0H U312 ( .A(n401), .B(n181), .Z(n183) );
  AO17SVTX1 U313 ( .A(m1[0]), .B(n175), .C(n515), .D(n174), .Z(n177) );
  AO1CDSVTX1 U314 ( .A(n139), .B(n138), .C(m1[6]), .D(m1[7]), .Z(n140) );
  ND3SVTX1 U315 ( .A(n137), .B(n515), .C(m1[2]), .Z(n138) );
  ND3SVTX1 U316 ( .A(n324), .B(m1[15]), .C(n82), .Z(n83) );
  NR3SVTX1 U317 ( .A(m1[8]), .B(m1[11]), .C(n95), .Z(n53) );
  F_ND2SVTX0H U318 ( .A(n49), .B(n82), .Z(n50) );
  ND3SVTX1 U319 ( .A(n515), .B(n175), .C(n174), .Z(n41) );
  NR3SVTX1 U320 ( .A(m1[7]), .B(m1[5]), .C(m1[4]), .Z(n20) );
  IVSVTX0H U321 ( .A(n21), .Z(n23) );
  ND3SVTX1 U322 ( .A(n193), .B(n167), .C(n144), .Z(n25) );
  AO7SVTX1 U323 ( .A(n249), .B(n109), .C(n123), .Z(n110) );
  B_ND2SVTX0H U324 ( .A(n108), .B(n107), .Z(n109) );
  NR2ASVTX1 U325 ( .A(m1[22]), .B(n111), .Z(n117) );
  AO20SVTX1 U326 ( .A(n456), .B(n200), .C(n199), .D(n198), .Z(n202) );
  AO20SVTX1 U327 ( .A(n170), .B(n184), .C(n169), .D(n168), .Z(n171) );
  AO20SVTX1 U328 ( .A(n225), .B(n224), .C(n223), .D(n294), .Z(n234) );
  IVSVTX0H U329 ( .A(m1[11]), .Z(n159) );
  IVSVTX2 U330 ( .A(n304), .Z(n218) );
  AO3SVTX1 U331 ( .A(n155), .B(n330), .C(n357), .D(n154), .Z(n332) );
  NR2SVTX0H U332 ( .A(n271), .B(n356), .Z(n257) );
  IVSVTX2 U333 ( .A(m1[17]), .Z(n132) );
  F_ND2SVTX0H U334 ( .A(n265), .B(n281), .Z(n210) );
  AO20SVTX1 U335 ( .A(n256), .B(n225), .C(n190), .D(n59), .Z(n61) );
  F_ND2SVTX0H U336 ( .A(n465), .B(n471), .Z(n466) );
  NR2SVTX0H U337 ( .A(m1[5]), .B(n467), .Z(n457) );
  NR2SVTX0H U338 ( .A(m1[7]), .B(n460), .Z(n461) );
  NR2SVTX0H U339 ( .A(m1[7]), .B(n538), .Z(n539) );
  F_ND2SVTX0H U340 ( .A(n536), .B(n535), .Z(n537) );
  NR2SVTX0H U341 ( .A(n534), .B(n538), .Z(n530) );
  F_ND2SVTX0H U342 ( .A(n129), .B(n454), .Z(n70) );
  ND2SVTX2 U343 ( .A(n159), .B(n449), .Z(n444) );
  ND4SVTX1 U344 ( .A(n501), .B(n500), .C(n499), .D(n498), .Z(n502) );
  AO11NSVTX2 U345 ( .A(n543), .B(n404), .C(n719), .D(n403), .E(n540), .F(
        m1[13]), .Z(n427) );
  FA1SVTX1 U346 ( .A(m1[20]), .B(n347), .CI(n346), .CO(n592), .Z(n589) );
  AO11NSVTX1 U347 ( .A(n388), .B(n244), .C(n719), .D(n243), .E(n540), .F(n401), 
        .Z(n347) );
  OR4SVTX1 U348 ( .A(n713), .B(n490), .C(n319), .D(n384), .Z(n346) );
  ND4SVTX1 U349 ( .A(n727), .B(n726), .C(n725), .D(n724), .Z(n734) );
  AO7SVTX2 U350 ( .A(n613), .B(n756), .C(n612), .Z(n620) );
  EOSVTX1 U351 ( .A(n653), .B(n652), .Z(m2[12]) );
  EOSVTX1 U352 ( .A(n757), .B(n756), .Z(m2[13]) );
  EOSVTX1 U353 ( .A(n661), .B(n660), .Z(m2[14]) );
  ENSVTX1 U354 ( .A(n621), .B(n620), .Z(m2[15]) );
  EOSVTX1 U355 ( .A(n642), .B(n641), .Z(m2[18]) );
  EOSVTX1 U356 ( .A(n637), .B(n636), .Z(m2[19]) );
  EOSVTX1 U357 ( .A(n628), .B(n627), .Z(m2[20]) );
  AO6SVTX1 U358 ( .A(n663), .B(n626), .C(n625), .Z(n627) );
  ND2SVTX4 U359 ( .A(n781), .B(n780), .Z(n782) );
  IVSVTX4 U360 ( .A(n487), .Z(n388) );
  IVSVTX2 U361 ( .A(m1[8]), .Z(n179) );
  IVSVTX2 U362 ( .A(m1[12]), .Z(n81) );
  IVSVTX2 U363 ( .A(m1[14]), .Z(n75) );
  F_ND2ASVTX2 U364 ( .A(m1[13]), .B(n75), .Z(n82) );
  IVSVTX2 U365 ( .A(n82), .Z(n167) );
  ND2SVTX4 U366 ( .A(n81), .B(n167), .Z(n21) );
  NR2SVTX2 U367 ( .A(m1[7]), .B(m1[6]), .Z(n199) );
  F_ND2ASVTX2 U368 ( .A(m1[11]), .B(n134), .Z(n49) );
  NR2SVTX2 U369 ( .A(n49), .B(n142), .Z(n3) );
  IVSVTX0H U370 ( .A(m1[2]), .Z(n488) );
  IVSVTX0H U371 ( .A(m1[0]), .Z(n2) );
  F_ND2ASVTX2 U372 ( .A(m1[1]), .B(n2), .Z(n137) );
  IVSVTX2 U373 ( .A(m1[3]), .Z(n476) );
  IVSVTX2 U374 ( .A(n476), .Z(n515) );
  ND4SVTX2 U375 ( .A(n3), .B(n184), .C(n488), .D(n6), .Z(n4) );
  NR2SVTX2 U376 ( .A(m1[23]), .B(m1[20]), .Z(n206) );
  NR2SVTX2 U377 ( .A(m1[19]), .B(m1[18]), .Z(n354) );
  IVSVTX4 U378 ( .A(n132), .Z(n324) );
  NR2SVTX2 U379 ( .A(n324), .B(m1[16]), .Z(n144) );
  ND2SVTX4 U380 ( .A(n354), .B(n144), .Z(n265) );
  NR2SVTX2 U381 ( .A(n265), .B(n285), .Z(n150) );
  ND2SVTX2 U382 ( .A(n206), .B(n150), .Z(n215) );
  NR2SVTX2 U383 ( .A(m1[12]), .B(m1[13]), .Z(n136) );
  F_ND2ASVTX2 U384 ( .A(m1[9]), .B(n134), .Z(n163) );
  IVSVTX2 U385 ( .A(m1[4]), .Z(n456) );
  AO7SVTX1 U386 ( .A(m1[2]), .B(n515), .C(m1[5]), .Z(n200) );
  ND2SVTX2 U387 ( .A(n136), .B(n9), .Z(n17) );
  IVSVTX0H U388 ( .A(m1[26]), .Z(n32) );
  AO7SVTX1 U389 ( .A(m1[15]), .B(n17), .C(n10), .Z(n63) );
  F_AN2SVTX2 U390 ( .A(n324), .B(m1[16]), .Z(n201) );
  IVSVTX0H U391 ( .A(n201), .Z(n11) );
  NR2ASVTX1 U392 ( .A(m1[23]), .B(n106), .Z(n209) );
  AO6SVTX2 U393 ( .A(n281), .B(n15), .C(n209), .Z(n64) );
  IVSVTX2 U394 ( .A(n352), .Z(n255) );
  AO7SVTX1 U395 ( .A(m1[1]), .B(m1[2]), .C(n515), .Z(n166) );
  IVSVTX0H U396 ( .A(n49), .Z(n193) );
  AO21SVTX1 U397 ( .A(m1[15]), .B(n324), .C(m1[16]), .D(n401), .Z(n22) );
  AO1SVTX1 U398 ( .A(n144), .B(n23), .C(n314), .D(n22), .Z(n24) );
  IVSVTX2 U399 ( .A(m1[19]), .Z(n168) );
  IVSVTX0H U400 ( .A(m1[25]), .Z(n775) );
  IVSVTX4 U401 ( .A(m1[22]), .Z(n330) );
  ND3SVTX2 U402 ( .A(n775), .B(n330), .C(n105), .Z(n190) );
  F_AN2SVTX2 U403 ( .A(m1[21]), .B(m1[20]), .Z(n38) );
  AO1ABSVTX1 U404 ( .A(n314), .B(n168), .C(n190), .D(n38), .Z(n27) );
  AO17SVTX2 U405 ( .A(n28), .B(n27), .C(n32), .D(n108), .Z(n66) );
  NR4SVTX2 U406 ( .A(m1[24]), .B(n32), .C(n123), .D(n31), .Z(n35) );
  IVSVTX0H U407 ( .A(n215), .Z(n33) );
  F_ND3SVTX2 U408 ( .A(n35), .B(n34), .C(n304), .Z(n410) );
  AO6SVTX1 U409 ( .A(n65), .B(n330), .C(n352), .Z(n58) );
  NR2SVTX2 U410 ( .A(n75), .B(n136), .Z(n92) );
  IVSVTX0H U411 ( .A(n92), .Z(n36) );
  AO7SVTX1 U412 ( .A(n184), .B(n36), .C(n170), .Z(n37) );
  ND4SVTX1 U413 ( .A(n324), .B(m1[26]), .C(n401), .D(n37), .Z(n45) );
  IVSVTX2 U414 ( .A(n38), .Z(n356) );
  IVSVTX0H U415 ( .A(m1[1]), .Z(n39) );
  AO6SVTX1 U416 ( .A(n178), .B(n41), .C(n194), .Z(n43) );
  IVSVTX0H U417 ( .A(m1[13]), .Z(n130) );
  NR3SVTX2 U418 ( .A(n45), .B(n356), .C(n44), .Z(n68) );
  NR2SVTX2 U419 ( .A(n324), .B(n401), .Z(n169) );
  NR3SVTX2 U420 ( .A(n168), .B(n169), .C(n330), .Z(n59) );
  NR2SVTX2 U421 ( .A(m1[25]), .B(n90), .Z(n219) );
  IVSVTX0H U422 ( .A(n219), .Z(n47) );
  ND3SVTX2 U423 ( .A(n295), .B(n327), .C(n46), .Z(n153) );
  IVSVTX0H U424 ( .A(n176), .Z(n95) );
  IVSVTX0H U425 ( .A(m1[6]), .Z(n48) );
  IVSVTX0H U426 ( .A(n77), .Z(n52) );
  AO3SVTX1 U427 ( .A(n76), .B(n515), .C(m1[4]), .D(m1[7]), .Z(n51) );
  AO8SVTX1 U428 ( .A(n53), .B(n52), .C(n51), .D(n50), .Z(n55) );
  AN4SVTX1 U429 ( .A(m1[16]), .B(m1[19]), .C(m1[22]), .D(m1[26]), .Z(n54) );
  AO7SVTX1 U430 ( .A(n56), .B(n55), .C(n54), .Z(n60) );
  F_ND2ASVTX2 U431 ( .A(m1[21]), .B(n149), .Z(n225) );
  AO7SVTX1 U432 ( .A(n352), .B(n61), .C(n60), .Z(n62) );
  ND4SVTX2 U433 ( .A(n64), .B(n219), .C(n63), .D(n62), .Z(n373) );
  ND4SVTX1 U434 ( .A(n119), .B(n105), .C(n330), .D(n65), .Z(n67) );
  ND3ABSVTX2 U435 ( .A(n68), .B(n67), .C(n66), .Z(n495) );
  IVSVTX0H U436 ( .A(m1[12]), .Z(n71) );
  NR2SVTX2 U437 ( .A(m1[9]), .B(n534), .Z(n129) );
  NR2SVTX2 U438 ( .A(m1[6]), .B(m1[5]), .Z(n454) );
  NR2SVTX2 U439 ( .A(n453), .B(n70), .Z(n529) );
  NR2SVTX2 U440 ( .A(m1[11]), .B(n524), .Z(n448) );
  NR2SVTX2 U441 ( .A(m1[15]), .B(n433), .Z(n428) );
  NR2SVTX2 U442 ( .A(n324), .B(n423), .Z(n400) );
  NR2SVTX2 U443 ( .A(m1[19]), .B(n389), .Z(n377) );
  NR2SVTX2 U444 ( .A(m1[21]), .B(n348), .Z(n322) );
  NR2SVTX2 U445 ( .A(m1[23]), .B(n241), .Z(n235) );
  ENSVTX0H U446 ( .A(m1[24]), .B(n235), .Z(n208) );
  F_ND2ASVTX2 U447 ( .A(n330), .B(n297), .Z(n73) );
  NR2ASVTX2 U448 ( .A(m1[22]), .B(n271), .Z(n74) );
  NR2SVTX2 U449 ( .A(n74), .B(n153), .Z(n102) );
  IVSVTX2 U450 ( .A(n102), .Z(n254) );
  ND4SVTX1 U451 ( .A(n515), .B(m1[5]), .C(m1[7]), .D(n76), .Z(n80) );
  AO7SVTX1 U452 ( .A(m1[6]), .B(m1[4]), .C(n77), .Z(n79) );
  AO8SVTX1 U453 ( .A(n80), .B(n179), .C(n79), .D(n78), .Z(n85) );
  AO1ABSVTX1 U454 ( .A(m1[14]), .B(n187), .C(n83), .D(n115), .Z(n84) );
  AO7SVTX2 U455 ( .A(n86), .B(n85), .C(n84), .Z(n88) );
  AO7SVTX1 U456 ( .A(n401), .B(n201), .C(n123), .Z(n87) );
  AO17SVTX2 U457 ( .A(n124), .B(n248), .C(n119), .D(n89), .Z(n112) );
  ND4ABCSVTX2 U458 ( .A(n258), .B(n90), .C(n254), .D(n112), .Z(n405) );
  IVSVTX0H U459 ( .A(n115), .Z(n91) );
  ND4SVTX1 U460 ( .A(n105), .B(n108), .C(n327), .D(n91), .Z(n104) );
  IVSVTX0H U461 ( .A(n96), .Z(n94) );
  AO21SVTX1 U462 ( .A(n95), .B(n94), .C(n93), .D(n92), .Z(n99) );
  ND4SVTX1 U463 ( .A(n96), .B(n160), .C(n176), .D(n465), .Z(n97) );
  AO20SVTX2 U464 ( .A(n515), .B(n175), .C(m1[4]), .D(n97), .Z(n98) );
  NR4ABSVTX1 U465 ( .A(m1[16]), .B(n401), .C(n115), .D(n149), .Z(n100) );
  IVSVTX0H U466 ( .A(n117), .Z(n103) );
  F_AO2SVTX1 U467 ( .A(n102), .B(n311), .C(n295), .D(n330), .Z(n362) );
  ND4ABSVTX2 U468 ( .A(n116), .B(n104), .C(n103), .D(n362), .Z(n341) );
  IVSVTX0H U469 ( .A(n116), .Z(n107) );
  NR2ASVTX2 U470 ( .A(n113), .B(n112), .Z(n369) );
  AO20SVTX2 U471 ( .A(n311), .B(n115), .C(n114), .D(n113), .Z(n406) );
  AO20SVTX1 U472 ( .A(m1[21]), .B(n116), .C(m1[22]), .D(n256), .Z(n118) );
  AO6ABSVTX1 U473 ( .A(n119), .B(n118), .C(n117), .Z(n125) );
  NR2ASVTX1 U474 ( .A(m1[23]), .B(n314), .Z(n211) );
  ND2SVTX2 U475 ( .A(n211), .B(n121), .Z(n122) );
  AO17CSVTX2 U476 ( .A(n124), .B(n213), .C(n123), .D(n122), .Z(n126) );
  NR2SVTX2 U477 ( .A(n125), .B(n126), .Z(n335) );
  NR2SVTX2 U478 ( .A(n406), .B(n335), .Z(n497) );
  IVSVTX4 U479 ( .A(n708), .Z(n489) );
  IVSVTX0H U480 ( .A(m1[15]), .Z(n131) );
  IVSVTX0H U481 ( .A(m1[2]), .Z(n475) );
  NR2SVTX2 U482 ( .A(m1[12]), .B(n444), .Z(n439) );
  ND2SVTX2 U483 ( .A(n130), .B(n439), .Z(n434) );
  NR2SVTX2 U484 ( .A(m1[14]), .B(n434), .Z(n429) );
  ND2SVTX2 U485 ( .A(n131), .B(n429), .Z(n424) );
  NR2SVTX2 U486 ( .A(m1[16]), .B(n424), .Z(n402) );
  NR2SVTX2 U487 ( .A(m1[20]), .B(n349), .Z(n323) );
  ND2SVTX2 U488 ( .A(n314), .B(n323), .Z(n242) );
  NR2SVTX2 U489 ( .A(m1[22]), .B(n242), .Z(n236) );
  ENSVTX0H U490 ( .A(m1[23]), .B(n236), .Z(n207) );
  IVSVTX0H U491 ( .A(n136), .Z(n141) );
  NR3SVTX2 U492 ( .A(n142), .B(n141), .C(n140), .Z(n145) );
  AO4SVTX2 U493 ( .A(n146), .B(n145), .C(n144), .D(n143), .Z(n282) );
  NR2ASVTX1 U494 ( .A(m1[23]), .B(n330), .Z(n148) );
  AO6CSVTX2 U495 ( .A(n155), .B(n268), .C(n148), .Z(n262) );
  IVSVTX0H U496 ( .A(n148), .Z(n222) );
  ND4SVTX1 U497 ( .A(n268), .B(n155), .C(n222), .D(n357), .Z(n152) );
  NR2ASVTX1 U498 ( .A(m1[23]), .B(n311), .Z(n151) );
  AO6CSVTX2 U499 ( .A(n150), .B(n149), .C(m1[23]), .Z(n228) );
  NR2SVTX2 U500 ( .A(n151), .B(n228), .Z(n221) );
  IVSVTX0H U501 ( .A(n153), .Z(n154) );
  NR2SVTX2 U502 ( .A(n332), .B(n156), .Z(n339) );
  NR2SVTX2 U503 ( .A(n157), .B(n255), .Z(n245) );
  IVSVTX0H U504 ( .A(n163), .Z(n161) );
  AO6SVTX1 U505 ( .A(n161), .B(n160), .C(n159), .Z(n162) );
  AO3SVTX1 U506 ( .A(m1[8]), .B(n163), .C(n162), .D(m1[12]), .Z(n164) );
  AO3SVTX2 U507 ( .A(n173), .B(n172), .C(n171), .D(m1[20]), .Z(n329) );
  AO8SVTX1 U508 ( .A(n179), .B(n178), .C(n177), .D(n176), .Z(n188) );
  NR2ASVTX1 U509 ( .A(m1[13]), .B(n183), .Z(n186) );
  AO6SVTX1 U510 ( .A(n201), .B(n401), .C(m1[19]), .Z(n182) );
  AO7SVTX1 U511 ( .A(n184), .B(n183), .C(n182), .Z(n185) );
  AO20SVTX2 U512 ( .A(n188), .B(n187), .C(n186), .D(n185), .Z(n278) );
  AO3SVTX2 U513 ( .A(n278), .B(n314), .C(n248), .D(n357), .Z(n364) );
  NR2ASVTX2 U514 ( .A(n189), .B(n364), .Z(n395) );
  IVSVTX0H U515 ( .A(n190), .Z(n353) );
  F_ND2SVTX0H U516 ( .A(m1[12]), .B(m1[13]), .Z(n195) );
  IVSVTX0H U517 ( .A(n191), .Z(n192) );
  AO7SVTX1 U518 ( .A(n193), .B(n195), .C(n192), .Z(n203) );
  IVSVTX0H U519 ( .A(n194), .Z(n197) );
  IVSVTX0H U520 ( .A(n195), .Z(n196) );
  AO7SVTX1 U521 ( .A(n203), .B(n202), .C(n201), .Z(n355) );
  NR2SVTX2 U522 ( .A(n256), .B(n273), .Z(n328) );
  AO7SVTX1 U523 ( .A(n354), .B(n272), .C(n328), .Z(n287) );
  AO17ASVTX2 U524 ( .A(n282), .B(n206), .C(n205), .D(n280), .Z(n491) );
  NR2SVTX2 U525 ( .A(n395), .B(n491), .Z(n382) );
  AO11NSVTX2 U526 ( .A(n543), .B(n208), .C(n719), .D(n207), .E(n540), .F(
        m1[19]), .Z(n321) );
  IVSVTX2 U527 ( .A(n252), .Z(n315) );
  NR2ASVTX1 U528 ( .A(n706), .B(n209), .Z(n261) );
  AO8SVTX1 U529 ( .A(n352), .B(n261), .C(n210), .D(n266), .Z(n229) );
  IVSVTX0H U530 ( .A(n229), .Z(n214) );
  F_AN2SVTX2 U531 ( .A(m1[25]), .B(n265), .Z(n298) );
  AO7SVTX1 U532 ( .A(n298), .B(n252), .C(n211), .Z(n212) );
  AO3SVTX1 U533 ( .A(n213), .B(n775), .C(n212), .D(n245), .Z(n232) );
  AO20SVTX2 U534 ( .A(n231), .B(n315), .C(n214), .D(n232), .Z(n371) );
  IVSVTX2 U535 ( .A(n245), .Z(n294) );
  AO7SVTX1 U536 ( .A(n255), .B(n215), .C(n294), .Z(n216) );
  AO7SVTX1 U537 ( .A(n315), .B(n706), .C(n216), .Z(n217) );
  AO17SVTX2 U538 ( .A(n219), .B(n218), .C(n352), .D(n217), .Z(n412) );
  ND4SVTX1 U539 ( .A(n245), .B(m1[25]), .C(n221), .D(n220), .Z(n485) );
  NR2ASVTX1 U540 ( .A(m1[23]), .B(n356), .Z(n227) );
  NR2ASVTX1 U541 ( .A(m1[25]), .B(n222), .Z(n223) );
  AO1SVTX1 U542 ( .A(n298), .B(n227), .C(n223), .D(n294), .Z(n233) );
  AO17ASVTX1 U543 ( .A(n315), .B(n227), .C(n226), .D(n234), .Z(n409) );
  F_AO2SVTX1 U544 ( .A(n228), .B(m1[25]), .C(m1[23]), .D(n252), .Z(n230) );
  AO1ABSVTX1 U545 ( .A(n311), .B(n231), .C(n230), .D(n229), .Z(n411) );
  AN3SVTX2 U546 ( .A(n309), .B(n233), .C(n232), .Z(n370) );
  AO20SVTX2 U547 ( .A(n304), .B(n255), .C(n294), .D(n234), .Z(n336) );
  NR3SVTX2 U548 ( .A(n411), .B(n370), .C(n336), .Z(n381) );
  ND4SVTX1 U549 ( .A(n412), .B(n485), .C(n409), .D(n381), .Z(n723) );
  ND3SVTX2 U550 ( .A(n405), .B(n383), .C(n497), .Z(n713) );
  EOSVTX0H U551 ( .A(m1[25]), .B(n715), .Z(n238) );
  OR2SVTX2 U552 ( .A(n240), .B(n239), .Z(n730) );
  EOSVTX0H U553 ( .A(m1[23]), .B(n241), .Z(n244) );
  EOSVTX2 U554 ( .A(m1[22]), .B(n242), .Z(n243) );
  IVSVTX0H U555 ( .A(n298), .Z(n246) );
  AO7SVTX1 U556 ( .A(n314), .B(n246), .C(n245), .Z(n247) );
  AO6ABSVTX1 U557 ( .A(n775), .B(n248), .C(n247), .Z(n313) );
  IVSVTX0H U558 ( .A(n249), .Z(n250) );
  NR2ASVTX1 U559 ( .A(m1[25]), .B(n250), .Z(n251) );
  AO1SVTX1 U560 ( .A(m1[20]), .B(n298), .C(n255), .D(n251), .Z(n303) );
  F_AO2SVTX1 U561 ( .A(n303), .B(n270), .C(m1[21]), .D(n297), .Z(n253) );
  AO21SVTX1 U562 ( .A(m1[24]), .B(n255), .C(n254), .D(n273), .Z(n306) );
  NR2SVTX2 U563 ( .A(n256), .B(n255), .Z(n267) );
  IVSVTX0H U564 ( .A(n267), .Z(n274) );
  AO21SVTX1 U565 ( .A(m1[22]), .B(n257), .C(n274), .D(n273), .Z(n310) );
  AO20SVTX2 U566 ( .A(n356), .B(n315), .C(n310), .D(n258), .Z(n259) );
  ND2SVTX2 U567 ( .A(n306), .B(n259), .Z(n722) );
  ND4SVTX2 U568 ( .A(n345), .B(n372), .C(n722), .D(n260), .Z(n490) );
  AO7SVTX1 U569 ( .A(n295), .B(n329), .C(n261), .Z(n264) );
  IVSVTX0H U570 ( .A(n262), .Z(n263) );
  ND3SVTX2 U571 ( .A(n357), .B(n264), .C(n263), .Z(n360) );
  AO7SVTX1 U572 ( .A(m1[21]), .B(n265), .C(m1[22]), .Z(n269) );
  NR2ASVTX1 U573 ( .A(m1[22]), .B(n270), .Z(n277) );
  AO3SVTX1 U574 ( .A(n305), .B(n277), .C(n292), .D(n276), .Z(n494) );
  NR2ASVTX1 U575 ( .A(n293), .B(n278), .Z(n279) );
  IVSVTX0H U576 ( .A(n280), .Z(n286) );
  AO6SVTX1 U577 ( .A(m1[23]), .B(n282), .C(n281), .Z(n284) );
  ND4SVTX1 U578 ( .A(n289), .B(n360), .C(n494), .D(n288), .Z(n319) );
  IVSVTX0H U579 ( .A(n290), .Z(n291) );
  IVSVTX0H U580 ( .A(n393), .Z(n318) );
  IVSVTX0H U581 ( .A(n292), .Z(n302) );
  NR2ASVTX1 U582 ( .A(n295), .B(n294), .Z(n300) );
  AO7SVTX1 U583 ( .A(n298), .B(n297), .C(n296), .Z(n299) );
  AO3SVTX2 U584 ( .A(n302), .B(n301), .C(n300), .D(n299), .Z(n419) );
  ND4SVTX1 U585 ( .A(m1[25]), .B(n309), .C(n304), .D(n303), .Z(n414) );
  IVSVTX0H U586 ( .A(n305), .Z(n308) );
  AO7SVTX1 U587 ( .A(n315), .B(n330), .C(n306), .Z(n307) );
  ND3SVTX2 U588 ( .A(n309), .B(n308), .C(n307), .Z(n340) );
  AO7SVTX1 U589 ( .A(n311), .B(n356), .C(n310), .Z(n312) );
  AO20SVTX2 U590 ( .A(n315), .B(n314), .C(n313), .D(n312), .Z(n368) );
  NR3ABSVTX2 U591 ( .A(n414), .B(n340), .C(n368), .Z(n726) );
  IVSVTX0H U592 ( .A(n316), .Z(n344) );
  ND4SVTX2 U593 ( .A(n318), .B(n495), .C(n419), .D(n317), .Z(n384) );
  ENSVTX0H U594 ( .A(m1[22]), .B(n322), .Z(n326) );
  ENSVTX0H U595 ( .A(m1[21]), .B(n323), .Z(n325) );
  AO11NSVTX1 U596 ( .A(n543), .B(n326), .C(n719), .D(n325), .E(n540), .F(n324), 
        .Z(n376) );
  AO3SVTX1 U597 ( .A(n330), .B(n329), .C(n328), .D(n327), .Z(n334) );
  IVSVTX0H U598 ( .A(n334), .Z(n331) );
  AN4SVTX1 U599 ( .A(n409), .B(n419), .C(n484), .D(n405), .Z(n500) );
  IVSVTX0H U600 ( .A(n335), .Z(n338) );
  IVSVTX0H U601 ( .A(n336), .Z(n337) );
  ND4SVTX1 U602 ( .A(n494), .B(n407), .C(n338), .D(n337), .Z(n343) );
  IVSVTX0H U603 ( .A(n339), .Z(n415) );
  ND4SVTX1 U604 ( .A(n500), .B(n345), .C(n722), .D(n396), .Z(n375) );
  NR2SVTX2 U605 ( .A(n590), .B(n589), .Z(n629) );
  EOSVTX0H U606 ( .A(m1[21]), .B(n348), .Z(n351) );
  EOSVTX0H U607 ( .A(m1[20]), .B(n349), .Z(n350) );
  AO3SVTX1 U608 ( .A(n354), .B(n356), .C(n353), .D(n352), .Z(n358) );
  IVSVTX0H U609 ( .A(n358), .Z(n365) );
  AO7SVTX1 U610 ( .A(n359), .B(n358), .C(n357), .Z(n361) );
  AO1SVTX1 U611 ( .A(n365), .B(n364), .C(n363), .D(n394), .Z(n501) );
  NR4ABSVTX1 U612 ( .A(n484), .B(n407), .C(n367), .D(n366), .Z(n374) );
  NR3SVTX2 U613 ( .A(n370), .B(n369), .C(n368), .Z(n397) );
  ND4SVTX1 U614 ( .A(n419), .B(n372), .C(n494), .D(n492), .Z(n721) );
  OR2SVTX2 U615 ( .A(n587), .B(n586), .Z(n638) );
  ENSVTX0H U616 ( .A(m1[20]), .B(n377), .Z(n380) );
  ENSVTX0H U617 ( .A(m1[19]), .B(n378), .Z(n379) );
  AO11NSVTX2 U618 ( .A(n543), .B(n380), .C(n719), .D(n379), .E(n540), .F(
        m1[15]), .Z(n399) );
  ND4SVTX1 U619 ( .A(n383), .B(n382), .C(n501), .D(n381), .Z(n385) );
  NR2SVTX2 U620 ( .A(n629), .B(n632), .Z(n626) );
  ND2SVTX2 U621 ( .A(n622), .B(n626), .Z(n595) );
  EOSVTX0H U622 ( .A(m1[19]), .B(n389), .Z(n392) );
  EOSVTX0H U623 ( .A(n401), .B(n390), .Z(n391) );
  NR2SVTX2 U624 ( .A(n577), .B(n576), .Z(n605) );
  ENSVTX0H U625 ( .A(n401), .B(n400), .Z(n404) );
  ENSVTX0H U626 ( .A(m1[17]), .B(n402), .Z(n403) );
  IVSVTX0H U627 ( .A(n406), .Z(n408) );
  ND4SVTX2 U628 ( .A(n410), .B(n409), .C(n408), .D(n407), .Z(n417) );
  ND4SVTX2 U629 ( .A(n415), .B(n492), .C(n414), .D(n413), .Z(n416) );
  ND3SVTX8 U630 ( .A(n420), .B(n419), .C(n483), .Z(n546) );
  NR2SVTX2 U631 ( .A(n575), .B(n574), .Z(n614) );
  NR2SVTX2 U632 ( .A(n605), .B(n614), .Z(n579) );
  EOSVTX0H U633 ( .A(m1[17]), .B(n423), .Z(n426) );
  EOSVTX0H U634 ( .A(m1[16]), .B(n424), .Z(n425) );
  AO11NSVTX2 U635 ( .A(n543), .B(n426), .C(n719), .D(n425), .E(n540), .F(
        m1[12]), .Z(n432) );
  NR2SVTX2 U636 ( .A(n573), .B(n572), .Z(n654) );
  ENSVTX0H U637 ( .A(m1[16]), .B(n428), .Z(n431) );
  ENSVTX0H U638 ( .A(m1[15]), .B(n429), .Z(n430) );
  AO11NSVTX2 U639 ( .A(n543), .B(n431), .C(n719), .D(n430), .E(n540), .F(
        m1[11]), .Z(n437) );
  F_FA1SVTX1 U640 ( .A(m1[14]), .B(n432), .CI(n546), .CO(n573), .Z(n570) );
  NR2SVTX2 U641 ( .A(n571), .B(n570), .Z(n657) );
  NR2SVTX2 U642 ( .A(n654), .B(n657), .Z(n608) );
  EOSVTX0H U643 ( .A(m1[15]), .B(n433), .Z(n436) );
  EOSVTX0H U644 ( .A(m1[14]), .B(n434), .Z(n435) );
  AO11NSVTX2 U645 ( .A(n543), .B(n436), .C(n719), .D(n435), .E(n540), .F(
        m1[10]), .Z(n442) );
  NR2SVTX2 U646 ( .A(n567), .B(n566), .Z(n643) );
  ENSVTX0H U647 ( .A(m1[14]), .B(n438), .Z(n441) );
  ENSVTX0H U648 ( .A(m1[13]), .B(n439), .Z(n440) );
  AO11NSVTX2 U649 ( .A(n543), .B(n441), .C(n719), .D(n440), .E(n540), .F(m1[9]), .Z(n447) );
  FA1SVTX1 U650 ( .A(m1[12]), .B(n442), .CI(n546), .CO(n567), .Z(n564) );
  NR2SVTX2 U651 ( .A(n565), .B(n564), .Z(n650) );
  NR2SVTX2 U652 ( .A(n643), .B(n650), .Z(n569) );
  EOSVTX0H U653 ( .A(m1[13]), .B(n443), .Z(n446) );
  EOSVTX0H U654 ( .A(m1[12]), .B(n444), .Z(n445) );
  AO11NSVTX2 U655 ( .A(n543), .B(n446), .C(n719), .D(n445), .E(n540), .F(m1[8]), .Z(n452) );
  F_FA1SVTX1 U656 ( .A(m1[11]), .B(n447), .CI(n546), .CO(n565), .Z(n562) );
  NR2SVTX2 U657 ( .A(n563), .B(n562), .Z(n669) );
  ENSVTX0H U658 ( .A(m1[12]), .B(n448), .Z(n451) );
  ENSVTX0H U659 ( .A(m1[11]), .B(n449), .Z(n450) );
  AO11NSVTX2 U660 ( .A(n543), .B(n451), .C(n708), .D(n450), .E(n540), .F(m1[7]), .Z(n528) );
  NR2SVTX2 U661 ( .A(n561), .B(n560), .Z(n674) );
  NR2SVTX2 U662 ( .A(n669), .B(n674), .Z(n646) );
  NR2SVTX2 U663 ( .A(n581), .B(n610), .Z(n583) );
  IVSVTX0H U664 ( .A(n453), .Z(n471) );
  IVSVTX0H U665 ( .A(n460), .Z(n535) );
  ENSVTX0H U666 ( .A(m1[7]), .B(n535), .Z(n459) );
  IVSVTX0H U667 ( .A(n455), .Z(n472) );
  ENSVTX0H U668 ( .A(m1[6]), .B(n457), .Z(n458) );
  AO11NSVTX2 U669 ( .A(n543), .B(n459), .C(n719), .D(n458), .E(n540), .F(m1[2]), .Z(n470) );
  ENSVTX0H U670 ( .A(m1[8]), .B(n461), .Z(n464) );
  IVSVTX0H U671 ( .A(n462), .Z(n538) );
  EOSVTX0H U672 ( .A(m1[7]), .B(n538), .Z(n463) );
  AO11NSVTX2 U673 ( .A(n543), .B(n464), .C(n719), .D(n463), .E(n540), .F(n515), 
        .Z(n545) );
  NR2SVTX2 U674 ( .A(n521), .B(n520), .Z(n696) );
  EOSVTX0H U675 ( .A(m1[6]), .B(n466), .Z(n469) );
  EOSVTX0H U676 ( .A(m1[5]), .B(n467), .Z(n468) );
  AO11NSVTX2 U677 ( .A(n543), .B(n469), .C(n719), .D(n468), .E(n540), .F(m1[1]), .Z(n514) );
  NR2SVTX2 U678 ( .A(n519), .B(n518), .Z(n758) );
  NR2SVTX2 U679 ( .A(n696), .B(n758), .Z(n523) );
  ENSVTX0H U680 ( .A(m1[5]), .B(n471), .Z(n474) );
  ENSVTX0H U681 ( .A(m1[4]), .B(n472), .Z(n473) );
  AO11NSVTX2 U682 ( .A(n543), .B(n474), .C(n719), .D(n473), .E(n540), .F(m1[0]), .Z(n510) );
  ENSVTX0H U683 ( .A(n475), .B(n515), .Z(n478) );
  ENSVTX0H U684 ( .A(n476), .B(m1[4]), .Z(n477) );
  AO2NSVTX1 U685 ( .A(n478), .B(n708), .C(n543), .D(n477), .Z(n486) );
  IVSVTX0H U686 ( .A(n479), .Z(n482) );
  OR2SVTX4 U687 ( .A(n510), .B(n509), .Z(n702) );
  ND3SVTX2 U688 ( .A(n485), .B(n484), .C(n483), .Z(n507) );
  HA1SVTX2 U689 ( .A(m1[1]), .B(n486), .CO(n513), .S(n506) );
  OR2SVTX2 U690 ( .A(n507), .B(n506), .Z(n768) );
  AO4SVTX1 U691 ( .A(n489), .B(n488), .C(n487), .D(n476), .Z(n505) );
  IVSVTX0H U692 ( .A(n490), .Z(n499) );
  IVSVTX0H U693 ( .A(n491), .Z(n493) );
  ND4SVTX1 U694 ( .A(n495), .B(n494), .C(n493), .D(n492), .Z(n496) );
  NR2ASVTX1 U695 ( .A(n497), .B(n496), .Z(n498) );
  OR2SVTX2 U696 ( .A(m1[0]), .B(n502), .Z(n504) );
  AO6NSVTX4 U697 ( .A(n768), .B(n771), .C(n508), .Z(n705) );
  FAS1SVTX2 U698 ( .A(m1[2]), .B(n513), .CI(n512), .CO(n517), .Z(n509) );
  F_FA1SVTX1 U699 ( .A(n515), .B(n514), .CI(n546), .CO(n519), .Z(n516) );
  NR2SVTX2 U700 ( .A(n517), .B(n516), .Z(n763) );
  EOSVTX0H U701 ( .A(m1[11]), .B(n524), .Z(n527) );
  EOSVTX0H U702 ( .A(m1[10]), .B(n525), .Z(n526) );
  AO11NSVTX2 U703 ( .A(n543), .B(n527), .C(n719), .D(n526), .E(n540), .F(m1[6]), .Z(n533) );
  FA1SVTX1 U704 ( .A(m1[9]), .B(n528), .CI(n546), .CO(n561), .Z(n554) );
  NR2SVTX2 U705 ( .A(n555), .B(n554), .Z(n677) );
  ENSVTX0H U706 ( .A(m1[10]), .B(n529), .Z(n532) );
  ENSVTX0H U707 ( .A(m1[9]), .B(n530), .Z(n531) );
  AO11NSVTX2 U708 ( .A(n543), .B(n532), .C(n708), .D(n531), .E(n540), .F(m1[5]), .Z(n544) );
  NR2SVTX2 U709 ( .A(n553), .B(n552), .Z(n682) );
  NR2SVTX2 U710 ( .A(n677), .B(n682), .Z(n557) );
  IVSVTX0H U711 ( .A(n534), .Z(n536) );
  EOSVTX0H U712 ( .A(m1[9]), .B(n537), .Z(n542) );
  ENSVTX0H U713 ( .A(m1[8]), .B(n539), .Z(n541) );
  AO11NSVTX2 U714 ( .A(n543), .B(n542), .C(n719), .D(n541), .E(n540), .F(m1[4]), .Z(n547) );
  F_FA1SVTX1 U715 ( .A(m1[6]), .B(n547), .CI(n546), .CO(n551), .Z(n548) );
  NR2SVTX2 U716 ( .A(n549), .B(n548), .Z(n688) );
  NR2SVTX2 U717 ( .A(n685), .B(n688), .Z(n603) );
  ND2SVTX2 U718 ( .A(n549), .B(n548), .Z(n693) );
  ND2SVTX2 U719 ( .A(n563), .B(n562), .Z(n671) );
  AO7SVTX2 U720 ( .A(n619), .B(n605), .C(n607), .Z(n578) );
  AO6SVTX2 U721 ( .A(n579), .B(n611), .C(n578), .Z(n580) );
  AO7SVTX4 U722 ( .A(n609), .B(n581), .C(n580), .Z(n582) );
  IVSVTX2 U723 ( .A(n639), .Z(n588) );
  AO6SVTX4 U724 ( .A(n638), .B(n640), .C(n588), .Z(n633) );
  ND2SVTX2 U725 ( .A(n590), .B(n589), .Z(n631) );
  AO6SVTX2 U726 ( .A(n625), .B(n622), .C(n593), .Z(n594) );
  IVSVTX0H U727 ( .A(n674), .Z(n597) );
  IVSVTX0H U728 ( .A(n682), .Z(n600) );
  IVSVTX2 U729 ( .A(n601), .Z(n694) );
  AO6SVTX2 U730 ( .A(n694), .B(n603), .C(n602), .Z(n681) );
  IVSVTX0H U731 ( .A(n605), .Z(n606) );
  IVSVTX0H U732 ( .A(n608), .Z(n613) );
  AO7SVTX2 U733 ( .A(n610), .B(n673), .C(n609), .Z(n659) );
  IVSVTX2 U734 ( .A(n659), .Z(n756) );
  IVSVTX0H U735 ( .A(n611), .Z(n612) );
  IVSVTX0H U736 ( .A(n619), .Z(n615) );
  IVSVTX2 U737 ( .A(n624), .Z(n663) );
  IVSVTX0H U738 ( .A(n629), .Z(n630) );
  IVSVTX0H U739 ( .A(n632), .Z(n635) );
  IVSVTX0H U740 ( .A(n633), .Z(n634) );
  AO6SVTX1 U741 ( .A(n663), .B(n635), .C(n634), .Z(n636) );
  AO6SVTX1 U742 ( .A(n663), .B(n1), .C(n640), .Z(n641) );
  IVSVTX0H U743 ( .A(n643), .Z(n644) );
  IVSVTX0H U744 ( .A(n646), .Z(n649) );
  IVSVTX0H U745 ( .A(n647), .Z(n648) );
  AO7SVTX2 U746 ( .A(n649), .B(n673), .C(n648), .Z(n667) );
  IVSVTX0H U747 ( .A(n666), .Z(n651) );
  AO6SVTX1 U748 ( .A(n667), .B(n665), .C(n651), .Z(n652) );
  IVSVTX0H U749 ( .A(n654), .Z(n655) );
  IVSVTX0H U750 ( .A(n755), .Z(n658) );
  AO6SVTX1 U751 ( .A(n659), .B(n754), .C(n658), .Z(n660) );
  ENSVTX0H U752 ( .A(n664), .B(n663), .Z(m2[17]) );
  ENSVTX0H U753 ( .A(n668), .B(n667), .Z(m2[11]) );
  IVSVTX0H U754 ( .A(n669), .Z(n670) );
  AO7SVTX1 U755 ( .A(n674), .B(n673), .C(n672), .Z(n675) );
  ENSVTX0H U756 ( .A(n676), .B(n675), .Z(m2[10]) );
  IVSVTX0H U757 ( .A(n677), .Z(n678) );
  AO7SVTX1 U758 ( .A(n682), .B(n681), .C(n680), .Z(n683) );
  ENSVTX0H U759 ( .A(n684), .B(n683), .Z(m2[8]) );
  IVSVTX0H U760 ( .A(n685), .Z(n686) );
  IVSVTX0H U761 ( .A(n688), .Z(n692) );
  IVSVTX0H U762 ( .A(n693), .Z(n689) );
  AO6SVTX1 U763 ( .A(n694), .B(n692), .C(n689), .Z(n690) );
  ENSVTX0H U764 ( .A(n695), .B(n694), .Z(m2[5]) );
  IVSVTX0H U765 ( .A(n696), .Z(n697) );
  AO7SVTX1 U766 ( .A(n758), .B(n761), .C(n760), .Z(n700) );
  ENSVTX0H U767 ( .A(n701), .B(n700), .Z(m2[4]) );
  ENSVTX0H U768 ( .A(n705), .B(n704), .Z(m2[1]) );
  AO7SVTX1 U769 ( .A(n776), .B(n706), .C(n774), .Z(n772) );
  NR2ASVTX1 U770 ( .A(m1[23]), .B(n776), .Z(n707) );
  OR3SVTX2 U771 ( .A(n708), .B(n388), .C(n707), .Z(n712) );
  IVSVTX0H U772 ( .A(n781), .Z(n743) );
  AO6NSVTX1 U773 ( .A(n717), .B(m1[22]), .C(n388), .Z(n737) );
  F_FA1SVTX1 U774 ( .A(m1[25]), .B(n712), .CI(n711), .CO(n709), .Z(n741) );
  NR2SVTX2 U775 ( .A(n742), .B(n741), .Z(n744) );
  IVSVTX0H U776 ( .A(n723), .Z(n724) );
  F_FA1SVTX1 U777 ( .A(m1[23]), .B(n735), .CI(n734), .CO(n739), .Z(n732) );
  F_FA1SVTX1 U778 ( .A(m1[24]), .B(n737), .CI(n736), .CO(n742), .Z(n738) );
  OR2SVTX2 U779 ( .A(n739), .B(n738), .Z(n784) );
  AO7SVTX8 U780 ( .A(n744), .B(n747), .C(n746), .Z(n780) );
  IVSVTX0H U781 ( .A(n744), .Z(n745) );
  IVSVTX0H U782 ( .A(n749), .Z(n750) );
  EOSVTX2 U783 ( .A(n753), .B(n752), .Z(m2[22]) );
  IVSVTX0H U784 ( .A(n758), .Z(n759) );
  IVSVTX0H U785 ( .A(n763), .Z(n764) );
  ENSVTX0H U786 ( .A(n771), .B(n770), .Z(m2[0]) );
  HA1SVTX1 U787 ( .A(m1[26]), .B(n772), .CO(n773), .S(n710) );
  IVSVTX0H U788 ( .A(n773), .Z(n779) );
  AO7SVTX1 U789 ( .A(n776), .B(n775), .C(n774), .Z(n777) );
  EOSVTX0H U790 ( .A(m1[27]), .B(n777), .Z(n778) );
endmodule


module remap_top ( num_i, rslt_o );
  input [31:0] num_i;
  output [31:0] rslt_o;
  wire   n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n374,
         n375, n377, n378, n379, n380;
  wire   [27:0] keyvalues_m1;

  remap re_map ( .m1(keyvalues_m1), .m2(rslt_o[26:0]) );
  AO3SVTX1 U198 ( .A(n319), .B(n366), .C(n307), .D(n306), .Z(keyvalues_m1[18])
         );
  MUX21NSVTX1 U199 ( .A(n315), .B(n304), .S(n378), .Z(n286) );
  IVSVTX0H U200 ( .A(n300), .Z(n273) );
  AO11NSVTX1 U201 ( .A(n310), .B(n348), .C(n311), .D(n229), .E(n285), .F(n371), 
        .Z(n304) );
  IVSVTX0H U202 ( .A(n269), .Z(n347) );
  MUX21NSVTX1 U203 ( .A(n321), .B(n320), .S(n378), .Z(n322) );
  IVSVTX0H U204 ( .A(n302), .Z(n316) );
  F_AO2SVTX1 U205 ( .A(n294), .B(num_i[6]), .C(rslt_o[28]), .D(n293), .Z(n326)
         );
  AO4SVTX1 U206 ( .A(n253), .B(n252), .C(n251), .D(n250), .Z(n289) );
  AO4SVTX1 U207 ( .A(n250), .B(n279), .C(n353), .D(n244), .Z(n254) );
  NR2ASVTX1 U208 ( .A(n355), .B(n351), .Z(n299) );
  IVSVTX2 U209 ( .A(n371), .Z(n323) );
  MUX21NSVTX1 U210 ( .A(n331), .B(n330), .S(rslt_o[28]), .Z(n333) );
  F_AO2SVTX1 U211 ( .A(n346), .B(n246), .C(n335), .D(n369), .Z(n247) );
  MUX21NSVTX1 U212 ( .A(n277), .B(n293), .S(n369), .Z(n332) );
  AO7SVTX1 U213 ( .A(n227), .B(n361), .C(n226), .Z(n372) );
  NR2ASVTX1 U214 ( .A(num_i[11]), .B(n361), .Z(n234) );
  IVSVTX4 U215 ( .A(n229), .Z(n292) );
  NR2SVTX4 U216 ( .A(rslt_o[29]), .B(rslt_o[28]), .Z(n371) );
  IVSVTX0H U217 ( .A(num_i[9]), .Z(n279) );
  NR2ASVTX4 U218 ( .A(rslt_o[29]), .B(rslt_o[28]), .Z(n229) );
  IVSVTX0H U219 ( .A(num_i[2]), .Z(n189) );
  OR2BSVTX4 U220 ( .A(n197), .B(n198), .Z(rslt_o[29]) );
  NR2ASVTX1 U221 ( .A(n194), .B(n259), .Z(n197) );
  NR2ASVTX2 U222 ( .A(n207), .B(n188), .Z(n204) );
  IVSVTX2 U223 ( .A(n353), .Z(n259) );
  IVSVTX0H U224 ( .A(num_i[11]), .Z(n218) );
  NR4SVTX2 U225 ( .A(num_i[4]), .B(num_i[7]), .C(num_i[5]), .D(num_i[6]), .Z(
        n207) );
  IVSVTX0H U226 ( .A(num_i[19]), .Z(n167) );
  IVSVTX0H U227 ( .A(n352), .Z(n364) );
  AO4SVTX1 U228 ( .A(n284), .B(n323), .C(n299), .D(n292), .Z(n230) );
  NR2ASVTX2 U229 ( .A(n259), .B(n298), .Z(n327) );
  F_AO2SVTX1 U230 ( .A(n294), .B(num_i[3]), .C(num_i[5]), .D(n327), .Z(n308)
         );
  IVSVTX4 U231 ( .A(rslt_o[27]), .Z(n378) );
  MUX21NSVTX2 U232 ( .A(n295), .B(n309), .S(n378), .Z(keyvalues_m1[4]) );
  AO3SVTX4 U233 ( .A(n319), .B(n292), .C(n291), .D(n290), .Z(keyvalues_m1[16])
         );
  F_ND2SVTX0H U234 ( .A(num_i[2]), .B(n204), .Z(n213) );
  B_ND2SVTX2 U235 ( .A(num_i[3]), .B(n204), .Z(n191) );
  ND2ASVTX4 U236 ( .A(rslt_o[31]), .B(rslt_o[30]), .Z(n361) );
  F_AO2SVTX1 U237 ( .A(rslt_o[30]), .B(num_i[16]), .C(num_i[8]), .D(n260), .Z(
        n282) );
  MUX21NSVTX1 U238 ( .A(n321), .B(n300), .S(rslt_o[27]), .Z(n301) );
  B_ND2SVTX2 U239 ( .A(n348), .B(n316), .Z(n290) );
  B_ND2SVTX1 U240 ( .A(n310), .B(n346), .Z(n271) );
  NR2ASVTX1 U241 ( .A(n374), .B(n298), .Z(n231) );
  MUX21NSVTX1 U242 ( .A(n237), .B(n312), .S(n245), .Z(n238) );
  AO1SVTX2 U243 ( .A(num_i[19]), .B(n253), .C(num_i[27]), .D(n234), .Z(n235)
         );
  B_ND2SVTX2 U244 ( .A(n233), .B(n232), .Z(n352) );
  AO17SVTX2 U245 ( .A(num_i[5]), .B(n227), .C(num_i[7]), .D(n206), .Z(n193) );
  IVSVTX2 U246 ( .A(n206), .Z(n188) );
  ND2ASVTX6 U247 ( .A(n225), .B(n253), .Z(rslt_o[30]) );
  AO6ASVTX2 U248 ( .A(n207), .B(n206), .C(n223), .Z(n198) );
  NR2ASVTX4 U249 ( .A(n224), .B(n223), .Z(n253) );
  B_ND2SVTX2 U250 ( .A(num_i[19]), .B(n200), .Z(n202) );
  NR4SVTX4 U251 ( .A(num_i[15]), .B(num_i[14]), .C(num_i[13]), .D(num_i[12]), 
        .Z(n196) );
  ND3SVTX2 U252 ( .A(n272), .B(n271), .C(n270), .Z(n300) );
  CTMUX21NSVTX4 U253 ( .A(n274), .B(n377), .S(rslt_o[27]), .Z(keyvalues_m1[24]) );
  AO7SVTX4 U254 ( .A(n324), .B(n366), .C(n286), .Z(keyvalues_m1[19]) );
  MUX21NSVTX1 U255 ( .A(n305), .B(n304), .S(rslt_o[27]), .Z(n307) );
  B_ND2SVTX2 U256 ( .A(n346), .B(n316), .Z(n317) );
  IVSVTX10 U257 ( .A(n215), .Z(rslt_o[28]) );
  ND3SVTX2 U258 ( .A(num_i[1]), .B(n189), .C(n204), .Z(n190) );
  IVSVTX2 U259 ( .A(n361), .Z(n343) );
  F_ND2ASVTX2 U260 ( .A(n353), .B(n198), .Z(n278) );
  IVSVTX2 U261 ( .A(num_i[10]), .Z(n251) );
  IVSVTX2 U262 ( .A(num_i[6]), .Z(n227) );
  MUX21NSVTX1 U263 ( .A(n315), .B(n320), .S(rslt_o[27]), .Z(n318) );
  MUX21NSVTX2 U264 ( .A(n380), .B(n370), .S(rslt_o[27]), .Z(keyvalues_m1[27])
         );
  AO1SVTX2 U265 ( .A(n346), .B(n372), .C(n231), .D(n230), .Z(n274) );
  MUX21NSVTX2 U266 ( .A(n337), .B(n338), .S(n378), .Z(keyvalues_m1[12]) );
  B_ND2SVTX2 U267 ( .A(n314), .B(n313), .Z(n320) );
  CTIVSVTX2 U268 ( .A(n267), .Z(n268) );
  AO7SVTX2 U269 ( .A(n282), .B(n298), .C(n247), .Z(n267) );
  B_ND2SVTX2 U270 ( .A(n289), .B(n378), .Z(n302) );
  CTIVSVTX2 U271 ( .A(n296), .Z(n284) );
  B_ND2SVTX2 U272 ( .A(n254), .B(rslt_o[27]), .Z(n319) );
  B_ND2SVTX2 U273 ( .A(n259), .B(rslt_o[29]), .Z(n280) );
  NR3SVTX2 U274 ( .A(n209), .B(n187), .C(n186), .Z(n192) );
  AO4SVTX2 U275 ( .A(n220), .B(n218), .C(n259), .D(n173), .Z(n209) );
  ND3SVTX2 U276 ( .A(n360), .B(n202), .C(n201), .Z(n203) );
  IVSVTX8 U277 ( .A(n170), .Z(n353) );
  F_ND2SVTX1 U278 ( .A(num_i[13]), .B(n362), .Z(n178) );
  B_ND2SVTX1 U279 ( .A(num_i[9]), .B(n251), .Z(n185) );
  NR4SVTX4 U280 ( .A(num_i[11]), .B(num_i[10]), .C(num_i[9]), .D(num_i[8]), 
        .Z(n221) );
  OR4ABCDSVTX8 U281 ( .A(n193), .B(n192), .C(n191), .D(n190), .Z(rslt_o[27])
         );
  CTMUX21NSVTX4 U282 ( .A(n332), .B(n325), .S(n378), .Z(keyvalues_m1[7]) );
  MUX22SVTX2 U283 ( .A(n334), .B(n333), .S(n378), .ZN(keyvalues_m1[9]) );
  NR2ASVTX6 U284 ( .A(n259), .B(n292), .Z(n294) );
  AO39SVTX2 U285 ( .A(n292), .B(n284), .C(n298), .D(n283), .E(n323), .F(n282), 
        .Z(n315) );
  AO7SVTX2 U286 ( .A(n220), .B(n251), .C(n205), .Z(n210) );
  NR2ASVTX6 U287 ( .A(n221), .B(n220), .Z(n206) );
  MUX21NSVTX4 U288 ( .A(n308), .B(n243), .S(n378), .Z(keyvalues_m1[2]) );
  AO2SVTX1 U289 ( .A(n260), .B(num_i[14]), .C(num_i[22]), .D(n259), .Z(n226)
         );
  CTMUX21NSVTX4 U290 ( .A(n337), .B(n268), .S(rslt_o[27]), .Z(keyvalues_m1[13]) );
  AO7SVTX2 U291 ( .A(n319), .B(n298), .C(n249), .Z(keyvalues_m1[14]) );
  AO11NSVTX1 U292 ( .A(n259), .B(num_i[20]), .C(n260), .D(num_i[12]), .E(
        num_i[4]), .F(n343), .Z(n296) );
  AO7SVTX2 U293 ( .A(n324), .B(n298), .C(n257), .Z(keyvalues_m1[15]) );
  CTMUX21NSVTX4 U294 ( .A(n274), .B(n273), .S(n378), .Z(keyvalues_m1[23]) );
  IVSVTX0H U295 ( .A(n265), .Z(n219) );
  AO4SVTX1 U296 ( .A(n245), .B(n217), .C(n279), .D(n278), .Z(n266) );
  F_ND2SVTX0H U297 ( .A(n229), .B(n316), .Z(n306) );
  AO7ABSVTX1 U298 ( .A(num_i[15]), .B(n259), .C(n248), .Z(n285) );
  F_ND2SVTX0H U299 ( .A(num_i[7]), .B(n260), .Z(n248) );
  AO2SVTX1 U300 ( .A(n260), .B(num_i[11]), .C(num_i[19]), .D(n259), .Z(n261)
         );
  AO7SVTX1 U301 ( .A(n345), .B(n361), .C(n240), .Z(n310) );
  AO2SVTX1 U302 ( .A(n260), .B(num_i[13]), .C(num_i[21]), .D(n259), .Z(n240)
         );
  F_AO2SVTX1 U303 ( .A(n294), .B(num_i[5]), .C(rslt_o[28]), .D(n281), .Z(n295)
         );
  F_MUX21NSVTX1 U304 ( .A(n266), .B(n330), .S(n369), .Z(n339) );
  AO7SVTX1 U305 ( .A(n299), .B(n298), .C(n297), .Z(n321) );
  AO4SVTX1 U306 ( .A(n361), .B(n264), .C(n236), .D(n250), .Z(n312) );
  AO6ABSVTX1 U307 ( .A(n279), .B(n361), .C(n242), .Z(n269) );
  F_AO2SVTX1 U308 ( .A(n294), .B(num_i[4]), .C(num_i[6]), .D(n327), .Z(n309)
         );
  NR2ASVTX1 U309 ( .A(n327), .B(n303), .Z(keyvalues_m1[1]) );
  F_ND2SVTX0H U310 ( .A(num_i[4]), .B(n327), .Z(n243) );
  MUX21NSVTX2 U311 ( .A(n326), .B(n295), .S(n378), .Z(keyvalues_m1[5]) );
  MUX21NSVTX2 U312 ( .A(n334), .B(n339), .S(rslt_o[27]), .Z(keyvalues_m1[10])
         );
  NR2ASVTX1 U313 ( .A(num_i[8]), .B(n361), .Z(n351) );
  IVSVTX4 U314 ( .A(n298), .Z(n348) );
  AO7SVTX1 U315 ( .A(n251), .B(n361), .C(n228), .Z(n374) );
  IVSVTX4 U316 ( .A(n346), .Z(n366) );
  B_ND2SVTX0H U317 ( .A(num_i[25]), .B(n179), .Z(n180) );
  ND3SVTX1 U318 ( .A(num_i[17]), .B(n252), .C(n200), .Z(n183) );
  AO6SVTX1 U319 ( .A(n353), .B(num_i[23]), .C(n177), .Z(n205) );
  AO17NSVTX2 U320 ( .A(n207), .B(num_i[3]), .C(num_i[7]), .D(n206), .Z(n208)
         );
  NR2ASVTX1 U321 ( .A(num_i[14]), .B(rslt_o[31]), .Z(n211) );
  AO2SVTX1 U322 ( .A(n200), .B(num_i[18]), .C(num_i[26]), .D(n199), .Z(n201)
         );
  IVSVTX2 U323 ( .A(num_i[22]), .Z(n182) );
  IVSVTX2 U324 ( .A(num_i[20]), .Z(n166) );
  NR2SVTX2 U325 ( .A(num_i[23]), .B(num_i[21]), .Z(n165) );
  ND3SVTX4 U326 ( .A(n182), .B(n166), .C(n165), .Z(n194) );
  IVSVTX2 U327 ( .A(num_i[18]), .Z(n252) );
  NR2SVTX2 U328 ( .A(num_i[17]), .B(num_i[16]), .Z(n172) );
  ND3SVTX2 U329 ( .A(n167), .B(n252), .C(n172), .Z(n174) );
  IVSVTX2 U330 ( .A(num_i[30]), .Z(n169) );
  IVSVTX2 U331 ( .A(num_i[29]), .Z(n340) );
  NR2SVTX2 U332 ( .A(num_i[31]), .B(num_i[28]), .Z(n168) );
  ND3SVTX4 U333 ( .A(n169), .B(n340), .C(n168), .Z(n195) );
  NR2SVTX2 U334 ( .A(num_i[27]), .B(num_i[26]), .Z(n179) );
  ND3ABSVTX4 U335 ( .A(num_i[24]), .B(num_i[25]), .C(n179), .Z(n222) );
  OR2SVTX4 U336 ( .A(n195), .B(n222), .Z(n170) );
  ND4ABSVTX8 U337 ( .A(n194), .B(n174), .C(n196), .D(n353), .Z(n220) );
  IVSVTX0H U338 ( .A(n194), .Z(n171) );
  ND4SVTX1 U339 ( .A(n172), .B(num_i[15]), .C(n252), .D(n171), .Z(n173) );
  NR3SVTX6 U340 ( .A(n195), .B(n222), .C(n194), .Z(n200) );
  ND2ASVTX8 U341 ( .A(n174), .B(n200), .Z(rslt_o[31]) );
  IVSVTX0H U342 ( .A(num_i[14]), .Z(n362) );
  IVSVTX0H U343 ( .A(num_i[27]), .Z(n176) );
  IVSVTX0H U344 ( .A(num_i[31]), .Z(n175) );
  AO7SVTX1 U345 ( .A(n176), .B(n195), .C(n175), .Z(n177) );
  AO3SVTX1 U346 ( .A(rslt_o[31]), .B(n178), .C(n202), .D(n205), .Z(n187) );
  AO4SVTX1 U347 ( .A(n195), .B(n180), .C(num_i[30]), .D(n340), .Z(n181) );
  AO8SVTX1 U348 ( .A(n353), .B(num_i[21]), .C(n182), .D(n181), .Z(n184) );
  AO3SVTX1 U349 ( .A(n185), .B(n220), .C(n184), .D(n183), .Z(n186) );
  IVSVTX2 U350 ( .A(n195), .Z(n199) );
  AO7SVTX4 U351 ( .A(n196), .B(rslt_o[31]), .C(n199), .Z(n223) );
  AO4SVTX1 U352 ( .A(n280), .B(n251), .C(n227), .D(n278), .Z(n277) );
  IVSVTX2 U353 ( .A(rslt_o[29]), .Z(n245) );
  AN2SVTX4 U354 ( .A(n353), .B(rslt_o[31]), .Z(n260) );
  AO2NSVTX1 U355 ( .A(num_i[4]), .B(n260), .C(num_i[12]), .D(n259), .Z(n246)
         );
  IVSVTX0H U356 ( .A(n246), .Z(n255) );
  IVSVTX0H U357 ( .A(num_i[8]), .Z(n276) );
  AO4SVTX1 U358 ( .A(n245), .B(n255), .C(n276), .D(n278), .Z(n336) );
  AO6SVTX1 U359 ( .A(n353), .B(num_i[22]), .C(num_i[30]), .Z(n360) );
  AO6SVTX1 U360 ( .A(n206), .B(num_i[6]), .C(n203), .Z(n214) );
  NR4SVTX2 U361 ( .A(n211), .B(n210), .C(n209), .D(n208), .Z(n212) );
  AN3SVTX4 U362 ( .A(n214), .B(n213), .C(n212), .Z(n215) );
  F_MUX21NSVTX1 U363 ( .A(n277), .B(n336), .S(rslt_o[28]), .Z(n334) );
  IVSVTX2 U364 ( .A(n260), .Z(n250) );
  IVSVTX0H U365 ( .A(num_i[5]), .Z(n345) );
  IVSVTX0H U366 ( .A(num_i[13]), .Z(n216) );
  AO4SVTX1 U367 ( .A(n250), .B(n345), .C(n353), .D(n216), .Z(n262) );
  IVSVTX0H U368 ( .A(n262), .Z(n217) );
  IVSVTX0H U369 ( .A(num_i[3]), .Z(n329) );
  AO4SVTX1 U370 ( .A(n250), .B(n329), .C(n353), .D(n218), .Z(n265) );
  IVSVTX0H U371 ( .A(num_i[7]), .Z(n264) );
  AO4SVTX1 U372 ( .A(n245), .B(n219), .C(n264), .D(n278), .Z(n330) );
  IVSVTX2 U373 ( .A(rslt_o[28]), .Z(n369) );
  AN2SVTX4 U374 ( .A(n245), .B(rslt_o[28]), .Z(n346) );
  NR2SVTX2 U375 ( .A(n221), .B(n220), .Z(n225) );
  IVSVTX0H U376 ( .A(n222), .Z(n224) );
  AO6SVTX1 U377 ( .A(n253), .B(num_i[18]), .C(num_i[26]), .Z(n228) );
  ND2SVTX4 U378 ( .A(rslt_o[29]), .B(rslt_o[28]), .Z(n298) );
  AO6SVTX1 U379 ( .A(n353), .B(num_i[16]), .C(num_i[24]), .Z(n355) );
  IVSVTX0H U380 ( .A(num_i[23]), .Z(n239) );
  IVSVTX0H U381 ( .A(rslt_o[31]), .Z(n233) );
  IVSVTX0H U382 ( .A(rslt_o[30]), .Z(n232) );
  AO7SVTX1 U383 ( .A(n329), .B(n352), .C(n235), .Z(n237) );
  IVSVTX0H U384 ( .A(num_i[15]), .Z(n236) );
  AO7SVTX2 U385 ( .A(n239), .B(n278), .C(n238), .Z(n350) );
  IVSVTX0H U386 ( .A(num_i[17]), .Z(n244) );
  IVSVTX0H U387 ( .A(num_i[25]), .Z(n241) );
  AO7SVTX1 U388 ( .A(n244), .B(rslt_o[30]), .C(n241), .Z(n242) );
  AO11SVTX2 U389 ( .A(n350), .B(rslt_o[28]), .C(n310), .D(n371), .E(n347), .F(
        n229), .Z(n377) );
  AO2ABSVTX1 U390 ( .C(num_i[6]), .D(n260), .A(n353), .B(n362), .Z(n258) );
  AO4SVTX1 U391 ( .A(n245), .B(n258), .C(n251), .D(n278), .Z(n335) );
  AO11NSVTX2 U392 ( .A(n285), .B(n229), .C(n262), .D(n346), .E(n265), .F(n371), 
        .Z(n256) );
  MUX21NSVTX2 U393 ( .A(n267), .B(n256), .S(rslt_o[27]), .Z(n249) );
  MUX21NSVTX2 U394 ( .A(n254), .B(n289), .S(rslt_o[27]), .Z(n324) );
  AO39SVTX1 U395 ( .A(n292), .B(n282), .C(n366), .D(n258), .E(n323), .F(n255), 
        .Z(n287) );
  MUX21NSVTX2 U396 ( .A(n287), .B(n256), .S(n378), .Z(n257) );
  AO39SVTX2 U397 ( .A(n366), .B(n282), .C(n298), .D(n284), .E(n323), .F(n258), 
        .Z(n305) );
  AO7SVTX1 U398 ( .A(n329), .B(n361), .C(n261), .Z(n311) );
  AO11NSVTX1 U399 ( .A(n285), .B(n346), .C(n311), .D(n348), .E(n262), .F(n371), 
        .Z(n288) );
  MUX21NSVTX2 U400 ( .A(n305), .B(n288), .S(n378), .Z(n263) );
  AO7SVTX2 U401 ( .A(n324), .B(n292), .C(n263), .Z(keyvalues_m1[17]) );
  AO4SVTX1 U402 ( .A(n280), .B(n264), .C(n329), .D(n278), .Z(n281) );
  AO11SVTX2 U403 ( .A(n266), .B(n369), .C(n265), .D(n346), .E(n285), .F(n348), 
        .Z(n337) );
  F_AO2SVTX1 U404 ( .A(n229), .B(n312), .C(n371), .D(n311), .Z(n272) );
  AO2ABSVTX1 U405 ( .C(num_i[23]), .D(n294), .A(n298), .B(n269), .Z(n270) );
  IVSVTX0H U406 ( .A(num_i[4]), .Z(n275) );
  AO4SVTX1 U407 ( .A(n280), .B(n276), .C(n278), .D(n275), .Z(n293) );
  AO4SVTX1 U408 ( .A(n280), .B(n279), .C(n278), .D(n345), .Z(n331) );
  F_MUX21NSVTX1 U409 ( .A(n331), .B(n281), .S(n369), .Z(n325) );
  IVSVTX0H U410 ( .A(n372), .Z(n283) );
  F_MUX21NSVTX1 U411 ( .A(n288), .B(n287), .S(n378), .Z(n291) );
  AO2SVTX2 U412 ( .A(n296), .B(n346), .C(n229), .D(n372), .Z(n297) );
  AO7SVTX4 U413 ( .A(n302), .B(n323), .C(n301), .Z(keyvalues_m1[22]) );
  F_MUX21NSVTX0H U414 ( .A(num_i[3]), .B(num_i[4]), .S(rslt_o[27]), .Z(n303)
         );
  F_MUX21NSVTX1 U415 ( .A(n309), .B(n308), .S(n378), .Z(keyvalues_m1[3]) );
  F_AO2SVTX1 U416 ( .A(n346), .B(n311), .C(n229), .D(n310), .Z(n314) );
  F_AO2SVTX1 U417 ( .A(n327), .B(num_i[23]), .C(n348), .D(n312), .Z(n313) );
  AO3SVTX4 U418 ( .A(n323), .B(n319), .C(n318), .D(n317), .Z(keyvalues_m1[20])
         );
  AO7SVTX4 U419 ( .A(n324), .B(n323), .C(n322), .Z(keyvalues_m1[21]) );
  MUX21NSVTX2 U420 ( .A(n326), .B(n325), .S(rslt_o[27]), .Z(keyvalues_m1[6])
         );
  IVSVTX0H U421 ( .A(n327), .Z(n328) );
  NR3SVTX2 U422 ( .A(n378), .B(n329), .C(n328), .Z(keyvalues_m1[0]) );
  MUX21NSVTX2 U423 ( .A(n332), .B(n333), .S(rslt_o[27]), .Z(keyvalues_m1[8])
         );
  F_MUX21NSVTX1 U424 ( .A(n336), .B(n335), .S(rslt_o[28]), .Z(n338) );
  MUX21NSVTX2 U425 ( .A(n339), .B(n338), .S(rslt_o[27]), .Z(keyvalues_m1[11])
         );
  IVSVTX0H U426 ( .A(num_i[21]), .Z(n341) );
  AO7SVTX1 U427 ( .A(n341), .B(rslt_o[30]), .C(n340), .Z(n342) );
  AO6SVTX1 U428 ( .A(n343), .B(num_i[13]), .C(n342), .Z(n344) );
  AO7SVTX1 U429 ( .A(n352), .B(n345), .C(n344), .Z(n349) );
  AO11SVTX2 U430 ( .A(n350), .B(n369), .C(n349), .D(n348), .E(n347), .F(n346), 
        .Z(n380) );
  IVSVTX0H U431 ( .A(n351), .Z(n359) );
  AO6SVTX1 U432 ( .A(n353), .B(num_i[20]), .C(num_i[28]), .Z(n354) );
  AO7SVTX1 U433 ( .A(n355), .B(rslt_o[29]), .C(n354), .Z(n357) );
  NR2ASVTX1 U434 ( .A(num_i[12]), .B(n361), .Z(n356) );
  AO1SVTX1 U435 ( .A(num_i[4]), .B(n364), .C(n357), .D(n356), .Z(n358) );
  AO7SVTX1 U436 ( .A(rslt_o[29]), .B(n359), .C(n358), .Z(n375) );
  IVSVTX0H U437 ( .A(n374), .Z(n367) );
  AO7SVTX1 U438 ( .A(n362), .B(n361), .C(n360), .Z(n363) );
  AO6SVTX1 U439 ( .A(num_i[6]), .B(n364), .C(n363), .Z(n365) );
  AO7SVTX1 U440 ( .A(n367), .B(n366), .C(n365), .Z(n368) );
  AO6SVTX1 U441 ( .A(n369), .B(n375), .C(n368), .Z(n370) );
  AO11SVTX2 U442 ( .A(n375), .B(rslt_o[28]), .C(n374), .D(n229), .E(n372), .F(
        n371), .Z(n379) );
  CTMUX21NSVTX4 U443 ( .A(n377), .B(n379), .S(rslt_o[27]), .Z(keyvalues_m1[25]) );
  MUX21NSVTX2 U444 ( .A(n380), .B(n379), .S(n378), .Z(keyvalues_m1[26]) );
endmodule

