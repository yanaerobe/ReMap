
module m_rangemapping ( N, O );
  input [31:0] N;
  output [31:0] O;
  wire   n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860;

  NR3ABSVTX1 U296 ( .A(n718), .B(n716), .C(n720), .Z(n706) );
  IVSVTX0H U297 ( .A(n770), .Z(n850) );
  IVSVTX0H U298 ( .A(n774), .Z(n776) );
  AO7SVTX1 U299 ( .A(n775), .B(n805), .C(n774), .Z(n783) );
  IVSVTX0H U300 ( .A(n789), .Z(n775) );
  EOSVTX1 U301 ( .A(n816), .B(n815), .Z(n818) );
  AO2NSVTX1 U302 ( .A(n498), .B(n490), .C(n494), .D(n493), .Z(n772) );
  AO11NSVTX1 U303 ( .A(n778), .B(n793), .C(n494), .D(n655), .E(n498), .F(n493), 
        .Z(n779) );
  HA1SVTX1 U304 ( .A(n768), .B(n489), .CO(n490), .S(n493) );
  AO11NSVTX1 U305 ( .A(n773), .B(n659), .C(n658), .D(n657), .E(n656), .F(n655), 
        .Z(n785) );
  HA1SVTX1 U306 ( .A(n492), .B(n491), .CO(n489), .S(n655) );
  AO7SVTX1 U307 ( .A(n295), .B(n284), .C(n290), .Z(n778) );
  AO11NSVTX1 U308 ( .A(n651), .B(n659), .C(n658), .D(n638), .E(n656), .F(n646), 
        .Z(n643) );
  AO7SVTX1 U309 ( .A(n461), .B(n295), .C(n294), .Z(n773) );
  AO11NSVTX1 U310 ( .A(n644), .B(n659), .C(n658), .D(n542), .E(n656), .F(n639), 
        .Z(n636) );
  AO6NSVTX1 U311 ( .A(n481), .B(n354), .C(n350), .Z(n781) );
  AO6NSVTX1 U312 ( .A(n481), .B(n336), .C(n332), .Z(n799) );
  AO6SVTX4 U313 ( .A(n742), .B(n211), .C(n607), .Z(n739) );
  AO11NSVTX1 U314 ( .A(n616), .B(n793), .C(n494), .D(n603), .E(n656), .F(n611), 
        .Z(n608) );
  EOSVTX1 U315 ( .A(n641), .B(n541), .Z(n545) );
  AO11NSVTX1 U316 ( .A(n609), .B(n793), .C(n658), .D(n595), .E(n656), .F(n604), 
        .Z(n601) );
  AO11SVTX1 U317 ( .A(N[5]), .B(n321), .C(n422), .D(N[21]), .E(n423), .F(N[13]), .Z(n345) );
  IVSVTX2 U318 ( .A(n819), .Z(n498) );
  MUX21NSVTX1 U319 ( .A(n391), .B(n396), .S(O[28]), .Z(n606) );
  AO2SVTX1 U320 ( .A(n423), .B(N[7]), .C(n422), .D(N[15]), .Z(n433) );
  IVSVTX0H U321 ( .A(n451), .Z(n408) );
  IVSVTX2 U322 ( .A(n284), .Z(n461) );
  BFSVTX4 U323 ( .A(n284), .Z(O[27]) );
  BFSVTX2 U324 ( .A(n285), .Z(n422) );
  IVSVTX0H U325 ( .A(n257), .Z(n234) );
  AO6SVTX1 U326 ( .A(N[3]), .B(n267), .C(n230), .Z(n231) );
  NR4SVTX2 U327 ( .A(N[27]), .B(N[26]), .C(N[25]), .D(N[24]), .Z(n216) );
  IVSVTX0H U328 ( .A(n651), .Z(n484) );
  ND2SVTX1 U329 ( .A(n556), .B(n419), .Z(n420) );
  AN2SVTX1 U330 ( .A(n339), .B(n504), .Z(n340) );
  ND2SVTX1 U331 ( .A(n401), .B(n400), .Z(n562) );
  AN2SVTX1 U332 ( .A(n811), .B(n810), .Z(n517) );
  NR2SVTX1 U333 ( .A(n799), .B(n798), .Z(n664) );
  IVSVTX2 U334 ( .A(n319), .Z(n321) );
  AO11NSVTX1 U335 ( .A(n582), .B(n793), .C(n494), .D(n572), .E(n498), .F(n574), 
        .Z(n575) );
  NR2SVTX1 U336 ( .A(n613), .B(n566), .Z(n561) );
  AO7SVTX1 U337 ( .A(n397), .B(n319), .C(n286), .Z(n329) );
  AO6ABSVTX1 U338 ( .A(O[29]), .B(n291), .C(n279), .Z(n311) );
  IVSVTX1 U339 ( .A(n369), .Z(n363) );
  IVSVTX2 U340 ( .A(O[28]), .Z(n426) );
  IVSVTX1 U341 ( .A(n284), .Z(n481) );
  AO7ABSVTX1 U342 ( .A(n658), .B(n597), .C(n596), .Z(n598) );
  AO2ASVTX1 U343 ( .C(n464), .D(n341), .A(n302), .B(O[28]), .Z(n295) );
  ND2SVTX1 U344 ( .A(n609), .B(n608), .Z(n738) );
  IVSVTX0H U345 ( .A(n844), .Z(n642) );
  ND2SVTX1 U346 ( .A(N[26]), .B(n381), .Z(n240) );
  AO6SVTX4 U347 ( .A(n751), .B(n749), .C(n600), .Z(n747) );
  ND2SVTX1 U348 ( .A(n690), .B(n689), .Z(n691) );
  AO6ABSVTX2 U349 ( .A(n632), .B(n212), .C(n631), .Z(n633) );
  EOSVTX1 U350 ( .A(n637), .B(n544), .Z(n549) );
  OR2SVTX2 U351 ( .A(n773), .B(n499), .Z(n358) );
  ND2SVTX2 U352 ( .A(n357), .B(n495), .Z(n499) );
  AO6ABSVTX1 U353 ( .A(n481), .B(n325), .C(n324), .Z(n326) );
  NR4SVTX2 U354 ( .A(N[27]), .B(N[25]), .C(N[24]), .D(n241), .Z(n243) );
  FA1SVTX4 U355 ( .A(n215), .B(n848), .CI(n847), .CO(n849), .Z(O[24]) );
  FA1SVTX4 U356 ( .A(n857), .B(n856), .CI(n855), .CO(n847), .Z(O[23]) );
  FA1SVTX4 U357 ( .A(n854), .B(n853), .CI(n852), .CO(n855), .Z(O[22]) );
  FA1SVTX4 U358 ( .A(n860), .B(n859), .CI(n858), .CO(n852), .Z(O[21]) );
  FA1SVTX2 U359 ( .A(n839), .B(n838), .CI(n837), .CO(n840), .Z(O[19]) );
  AO6SVTX2 U360 ( .A(n689), .B(n692), .C(n674), .Z(n833) );
  IVSVTX1 U361 ( .A(n690), .Z(n674) );
  ND2SVTX2 U362 ( .A(n805), .B(n821), .Z(n774) );
  FA1SVTX1 U363 ( .A(n828), .B(n827), .CI(n826), .CO(n839), .Z(n685) );
  ND2SVTX2 U364 ( .A(n494), .B(n775), .Z(n792) );
  EOSVTX4 U365 ( .A(n492), .B(n661), .Z(n789) );
  NR2SVTX2 U366 ( .A(n492), .B(n661), .Z(n662) );
  ND2SVTX4 U367 ( .A(n800), .B(n801), .Z(n661) );
  AO7SVTX6 U368 ( .A(n812), .B(n815), .C(n814), .Z(n801) );
  ND2ASVTX6 U369 ( .A(n654), .B(n653), .Z(n682) );
  IVSVTX2 U370 ( .A(n681), .Z(n660) );
  AO6ABSVTX2 U371 ( .A(n481), .B(n480), .C(n479), .Z(n482) );
  ND3ABSVTX4 U372 ( .A(n272), .B(n271), .C(n270), .Z(n284) );
  ND3SVTX2 U373 ( .A(N[17]), .B(n282), .C(n257), .Z(n258) );
  ND3SVTX2 U374 ( .A(N[1]), .B(n380), .C(n267), .Z(n268) );
  FA1SVTX4 U375 ( .A(n851), .B(n850), .CI(n849), .CO(n835), .Z(O[25]) );
  AO7SVTX2 U376 ( .A(n834), .B(n833), .C(n832), .Z(n837) );
  AN2SVTX2 U377 ( .A(n784), .B(n783), .Z(n215) );
  FA1SVTX2 U378 ( .A(n677), .B(n676), .CI(n675), .CO(n686), .Z(n692) );
  ND2SVTX2 U379 ( .A(n792), .B(n804), .Z(n770) );
  ND3ABSVTX4 U380 ( .A(n652), .B(n664), .C(n672), .Z(n653) );
  AO7SVTX6 U381 ( .A(n758), .B(n761), .C(n760), .Z(n672) );
  AO7SVTX6 U382 ( .A(n727), .B(n730), .C(n729), .Z(n725) );
  AO6SVTX6 U383 ( .A(n734), .B(n732), .C(n614), .Z(n730) );
  AO6SVTX2 U384 ( .A(n519), .B(n518), .C(n517), .Z(n667) );
  AO7SVTX4 U385 ( .A(n736), .B(n739), .C(n738), .Z(n734) );
  AO7SVTX2 U386 ( .A(n522), .B(n514), .C(n513), .Z(n519) );
  OR2SVTX2 U387 ( .A(n773), .B(n772), .Z(n800) );
  AO7SVTX6 U388 ( .A(n744), .B(n747), .C(n746), .Z(n742) );
  OR2SVTX2 U389 ( .A(n786), .B(n785), .Z(n680) );
  NR2SVTX2 U390 ( .A(n651), .B(n650), .Z(n758) );
  NR2SVTX2 U391 ( .A(n644), .B(n643), .Z(n763) );
  AO7SVTX4 U392 ( .A(n753), .B(n756), .C(n755), .Z(n751) );
  ENSVTX1 U393 ( .A(n811), .B(n511), .Z(n526) );
  EOSVTX2 U394 ( .A(n630), .B(n548), .Z(n552) );
  AO6SVTX4 U395 ( .A(n592), .B(n591), .C(n590), .Z(n756) );
  EOSVTX1 U396 ( .A(n628), .B(n551), .Z(n618) );
  AO7SVTX2 U397 ( .A(n585), .B(n584), .C(n583), .Z(n592) );
  AO6SVTX2 U398 ( .A(n213), .B(n580), .C(n579), .Z(n584) );
  OR2SVTX2 U399 ( .A(n507), .B(n358), .Z(n488) );
  AN2SVTX2 U400 ( .A(n576), .B(n575), .Z(n580) );
  ENSVTX1 U401 ( .A(n602), .B(n567), .Z(n586) );
  ND2SVTX1 U402 ( .A(n529), .B(n528), .Z(n530) );
  ND2SVTX2 U403 ( .A(n509), .B(n340), .Z(n507) );
  BFSVTX2 U404 ( .A(n494), .Z(n658) );
  IVSVTX2 U405 ( .A(n214), .Z(n659) );
  ND2SVTX1 U406 ( .A(n504), .B(n509), .Z(n505) );
  IVSVTX1 U407 ( .A(n644), .Z(n463) );
  OR2SVTX2 U408 ( .A(n822), .B(n678), .Z(n214) );
  ND2SVTX1 U409 ( .A(n392), .B(n564), .Z(n393) );
  IVSVTX2 U410 ( .A(n778), .Z(n492) );
  ND2SVTX2 U411 ( .A(n550), .B(n432), .Z(n546) );
  IVSVTX2 U412 ( .A(n625), .Z(n550) );
  AO7SVTX2 U413 ( .A(n439), .B(O[27]), .C(n438), .Z(n630) );
  ND2SVTX1 U414 ( .A(n361), .B(n360), .Z(n367) );
  AO6ABSVTX2 U415 ( .A(n481), .B(n472), .C(n471), .Z(n473) );
  AO4SVTX2 U416 ( .A(n375), .B(n364), .C(n376), .D(n363), .Z(n589) );
  NR2ASVTX2 U417 ( .A(n422), .B(n435), .Z(n384) );
  ND2SVTX1 U418 ( .A(N[4]), .B(n423), .Z(n412) );
  AO2SVTX2 U419 ( .A(n423), .B(N[1]), .C(n422), .D(N[9]), .Z(n440) );
  AN2BSVTX2 U420 ( .A(n226), .B(O[31]), .Z(n238) );
  AO6ASVTX2 U421 ( .A(n269), .B(n268), .C(O[31]), .Z(n271) );
  ND4ABCSVTX4 U422 ( .A(N[17]), .B(N[16]), .C(n218), .D(n257), .Z(O[31]) );
  NR2SVTX2 U423 ( .A(n217), .B(n422), .Z(n221) );
  NR2ASVTX4 U424 ( .A(n217), .B(n285), .Z(n257) );
  NR2SVTX1 U425 ( .A(N[10]), .B(n261), .Z(n263) );
  NR4SVTX4 U426 ( .A(N[11]), .B(N[10]), .C(N[9]), .D(N[8]), .Z(n239) );
  NR4SVTX6 U427 ( .A(N[30]), .B(N[31]), .C(N[29]), .D(N[28]), .Z(n381) );
  NR4SVTX6 U428 ( .A(N[14]), .B(N[15]), .C(N[13]), .D(N[12]), .Z(n264) );
  IVSVTX2 U429 ( .A(N[2]), .Z(n380) );
  AO4SVTX2 U430 ( .A(n319), .B(n406), .C(n404), .D(n248), .Z(n342) );
  AO2SVTX2 U431 ( .A(n423), .B(N[0]), .C(n422), .D(N[8]), .Z(n436) );
  AO11SVTX2 U432 ( .A(n448), .B(n468), .C(n429), .D(n466), .E(n474), .F(n464), 
        .Z(n439) );
  IVSVTX2 U433 ( .A(n662), .Z(n794) );
  AO1SVTX2 U434 ( .A(n407), .B(n342), .C(n253), .D(n252), .Z(n302) );
  AO20SVTX1 U435 ( .A(n403), .B(n298), .C(n251), .D(n407), .Z(n252) );
  AO7NSVTX1 U436 ( .A(n250), .B(O[30]), .C(n249), .Z(n251) );
  IVSVTX2 U437 ( .A(n423), .Z(n404) );
  AN2SVTX1 U438 ( .A(O[27]), .B(O[28]), .Z(n409) );
  ND2SVTX1 U439 ( .A(n466), .B(n341), .Z(n300) );
  AO11NSVTX1 U440 ( .A(n623), .B(n793), .C(n494), .D(n610), .E(n656), .F(n617), 
        .Z(n615) );
  AO11NSVTX1 U441 ( .A(n656), .B(n618), .C(n659), .D(n625), .E(n658), .F(n617), 
        .Z(n619) );
  AO11NSVTX1 U442 ( .A(n788), .B(n659), .C(n658), .D(n645), .E(n656), .F(n526), 
        .Z(n650) );
  AO7SVTX2 U443 ( .A(n817), .B(n679), .C(n663), .Z(n673) );
  ND2SVTX1 U444 ( .A(n814), .B(n813), .Z(n816) );
  NR2SVTX1 U445 ( .A(n616), .B(n615), .Z(n727) );
  ND2SVTX1 U446 ( .A(n616), .B(n615), .Z(n729) );
  ND2SVTX1 U447 ( .A(n620), .B(n619), .Z(n724) );
  OR2SVTX1 U448 ( .A(n620), .B(n619), .Z(n723) );
  ND2SVTX1 U449 ( .A(n651), .B(n650), .Z(n760) );
  NR2ASVTX2 U450 ( .A(n671), .B(n817), .Z(n675) );
  ND2SVTX1 U451 ( .A(n666), .B(n665), .Z(n670) );
  EOSVTX1 U452 ( .A(n784), .B(n783), .Z(n856) );
  IVSVTX0H U453 ( .A(n576), .Z(n360) );
  AO4SVTX2 U454 ( .A(n404), .B(n403), .C(n402), .D(n256), .Z(n451) );
  ND2SVTX1 U455 ( .A(n466), .B(n469), .Z(n328) );
  ND2SVTX1 U456 ( .A(n468), .B(n341), .Z(n344) );
  NR2ASVTX1 U457 ( .A(n362), .B(n363), .Z(n576) );
  ND2SVTX1 U458 ( .A(n556), .B(n555), .Z(n558) );
  AO4SVTX1 U459 ( .A(n440), .B(n407), .C(n394), .D(n405), .Z(n415) );
  NR2SVTX1 U460 ( .A(O[27]), .B(n426), .Z(n417) );
  IVSVTX0H U461 ( .A(N[5]), .Z(n394) );
  AO7SVTX2 U462 ( .A(n373), .B(n372), .C(n371), .Z(n594) );
  AO6CSVTX1 U463 ( .A(n672), .B(n668), .C(n667), .Z(n669) );
  ND2SVTX1 U464 ( .A(n681), .B(n680), .Z(n683) );
  AO6ABSVTX1 U465 ( .A(n284), .B(n349), .C(n293), .Z(n294) );
  NR2SVTX1 U466 ( .A(N[26]), .B(n254), .Z(n255) );
  FA1SVTX1 U467 ( .A(n831), .B(n830), .CI(n829), .CO(n842), .Z(n838) );
  AO7CSVTX1 U468 ( .A(n822), .B(n821), .C(n820), .Z(n829) );
  NR2SVTX1 U469 ( .A(n819), .B(n662), .Z(n820) );
  AO7SVTX1 U470 ( .A(n250), .B(n234), .C(n233), .Z(n235) );
  ND2SVTX1 U471 ( .A(N[22]), .B(n256), .Z(n228) );
  ND2SVTX1 U472 ( .A(N[18]), .B(n257), .Z(n227) );
  IVSVTX0H U473 ( .A(N[30]), .Z(n303) );
  ND2SVTX1 U474 ( .A(n738), .B(n737), .Z(n740) );
  ND2SVTX1 U475 ( .A(n733), .B(n732), .Z(n735) );
  ND2SVTX1 U476 ( .A(n729), .B(n728), .Z(n731) );
  ND2SVTX1 U477 ( .A(n724), .B(n723), .Z(n726) );
  ND2SVTX1 U478 ( .A(n719), .B(n718), .Z(n710) );
  ND2SVTX1 U479 ( .A(n717), .B(n716), .Z(n722) );
  ND2SVTX1 U480 ( .A(n704), .B(n703), .Z(n709) );
  ND2SVTX1 U481 ( .A(n699), .B(n698), .Z(n701) );
  ND2SVTX1 U482 ( .A(n765), .B(n764), .Z(n767) );
  ND2SVTX1 U483 ( .A(n694), .B(n693), .Z(n696) );
  ND2SVTX1 U484 ( .A(n760), .B(n759), .Z(n762) );
  ND2SVTX1 U485 ( .A(n832), .B(n687), .Z(n688) );
  OR2SVTX1 U486 ( .A(n606), .B(n605), .Z(n211) );
  AO7NSVTX1 U487 ( .A(n702), .B(n707), .C(n704), .Z(n212) );
  OR2SVTX2 U488 ( .A(n578), .B(n577), .Z(n213) );
  IVSVTX1 U489 ( .A(n553), .Z(n718) );
  NR2SVTX1 U490 ( .A(n623), .B(n622), .Z(n553) );
  NR4SVTX2 U491 ( .A(N[23]), .B(N[22]), .C(N[21]), .D(N[20]), .Z(n217) );
  ND2SVTX4 U492 ( .A(n216), .B(n381), .Z(n285) );
  NR4SVTX2 U493 ( .A(N[4]), .B(N[5]), .C(N[6]), .D(N[7]), .Z(n222) );
  ND2SVTX2 U494 ( .A(n239), .B(n264), .Z(n266) );
  IVSVTX2 U495 ( .A(N[19]), .Z(n250) );
  IVSVTX2 U496 ( .A(N[18]), .Z(n282) );
  ND2SVTX2 U497 ( .A(n250), .B(n282), .Z(n218) );
  NR3SVTX2 U498 ( .A(n222), .B(n266), .C(O[31]), .Z(n220) );
  IVSVTX0H U499 ( .A(n381), .Z(n219) );
  AO6ABSVTX2 U500 ( .A(n264), .B(O[31]), .C(n219), .Z(n242) );
  ND3ABSVTX4 U501 ( .A(n221), .B(n220), .C(n242), .Z(O[29]) );
  NR2ASVTX2 U502 ( .A(n222), .B(n266), .Z(n267) );
  IVSVTX0H U503 ( .A(n267), .Z(n225) );
  NR2ASVTX1 U504 ( .A(N[6]), .B(n266), .Z(n223) );
  AO1SVTX1 U505 ( .A(n264), .B(N[10]), .C(N[14]), .D(n223), .Z(n224) );
  AO7SVTX1 U506 ( .A(n380), .B(n225), .C(n224), .Z(n226) );
  IVSVTX0H U507 ( .A(n285), .Z(n256) );
  ND4SVTX2 U508 ( .A(n303), .B(n240), .C(n228), .D(n227), .Z(n237) );
  IVSVTX0H U509 ( .A(N[7]), .Z(n406) );
  AO6SVTX1 U510 ( .A(n264), .B(N[11]), .C(N[15]), .Z(n229) );
  AO7SVTX1 U511 ( .A(n406), .B(n266), .C(n229), .Z(n230) );
  NR2SVTX2 U512 ( .A(n231), .B(O[31]), .Z(n236) );
  NR2ASVTX1 U513 ( .A(N[23]), .B(n285), .Z(n232) );
  AO1SVTX1 U514 ( .A(n381), .B(N[27]), .C(N[31]), .D(n232), .Z(n233) );
  NR2SVTX2 U515 ( .A(n236), .B(n235), .Z(n270) );
  ND3ABSVTX6 U516 ( .A(n238), .B(n237), .C(n270), .Z(O[28]) );
  ND2SVTX4 U517 ( .A(O[29]), .B(n426), .Z(n435) );
  IVSVTX2 U518 ( .A(n435), .Z(n464) );
  IVSVTX0H U519 ( .A(N[1]), .Z(n374) );
  IVSVTX2 U520 ( .A(O[31]), .Z(n280) );
  IVSVTX0H U521 ( .A(n239), .Z(n244) );
  IVSVTX0H U522 ( .A(n240), .Z(n241) );
  AN2SVTX2 U523 ( .A(n243), .B(n242), .Z(n247) );
  AO7ABSVTX2 U524 ( .A(n280), .B(n244), .C(n247), .Z(O[30]) );
  NR2ASVTX2 U525 ( .A(n280), .B(O[30]), .Z(n307) );
  IVSVTX2 U526 ( .A(n307), .Z(n298) );
  IVSVTX0H U527 ( .A(O[30]), .Z(n296) );
  IVSVTX0H U528 ( .A(N[9]), .Z(n261) );
  IVSVTX0H U529 ( .A(N[25]), .Z(n254) );
  AO7SVTX1 U530 ( .A(n261), .B(O[31]), .C(n254), .Z(n245) );
  AO6SVTX1 U531 ( .A(n296), .B(N[17]), .C(n245), .Z(n246) );
  AO7SVTX2 U532 ( .A(n374), .B(n298), .C(n246), .Z(n341) );
  IVSVTX2 U533 ( .A(O[29]), .Z(n407) );
  ND2ASVTX2 U534 ( .A(O[31]), .B(O[30]), .Z(n319) );
  AN2SVTX4 U535 ( .A(O[31]), .B(n247), .Z(n423) );
  IVSVTX0H U536 ( .A(N[15]), .Z(n248) );
  ND2ASVTX2 U537 ( .A(O[29]), .B(n422), .Z(n405) );
  NR2ASVTX1 U538 ( .A(N[23]), .B(n405), .Z(n253) );
  IVSVTX0H U539 ( .A(N[3]), .Z(n403) );
  AO6SVTX1 U540 ( .A(n280), .B(N[11]), .C(N[27]), .Z(n249) );
  AO2SVTX1 U541 ( .A(n381), .B(n255), .C(N[29]), .D(n303), .Z(n260) );
  IVSVTX0H U542 ( .A(N[22]), .Z(n304) );
  ND3SVTX2 U543 ( .A(N[21]), .B(n304), .C(n256), .Z(n259) );
  ND3SVTX2 U544 ( .A(n260), .B(n259), .C(n258), .Z(n272) );
  IVSVTX0H U545 ( .A(N[14]), .Z(n262) );
  AO2SVTX1 U546 ( .A(n264), .B(n263), .C(N[13]), .D(n262), .Z(n265) );
  AO21SVTX1 U547 ( .A(N[6]), .B(n394), .C(n266), .D(n265), .Z(n269) );
  IVSVTX0H U548 ( .A(N[16]), .Z(n274) );
  AO6SVTX1 U549 ( .A(n280), .B(N[8]), .C(N[24]), .Z(n273) );
  AO7SVTX1 U550 ( .A(n274), .B(O[30]), .C(n273), .Z(n275) );
  AO6SVTX1 U551 ( .A(n307), .B(N[0]), .C(n275), .Z(n291) );
  IVSVTX0H U552 ( .A(N[12]), .Z(n278) );
  ND2SVTX2 U553 ( .A(N[4]), .B(n307), .Z(n277) );
  AO6SVTX1 U554 ( .A(n423), .B(N[20]), .C(N[28]), .Z(n276) );
  AO3SVTX1 U555 ( .A(n278), .B(n319), .C(n277), .D(n276), .Z(n279) );
  AO6SVTX1 U556 ( .A(n280), .B(N[10]), .C(N[26]), .Z(n281) );
  AO7SVTX1 U557 ( .A(n282), .B(O[30]), .C(n281), .Z(n283) );
  AO6SVTX1 U558 ( .A(N[2]), .B(n307), .C(n283), .Z(n309) );
  AO4SVTX1 U559 ( .A(n311), .B(n426), .C(n309), .D(n435), .Z(n313) );
  IVSVTX0H U560 ( .A(N[6]), .Z(n397) );
  AO2SVTX1 U561 ( .A(n423), .B(N[14]), .C(n422), .D(N[22]), .Z(n286) );
  IVSVTX0H U562 ( .A(n329), .Z(n288) );
  OR2SVTX2 U563 ( .A(O[29]), .B(O[28]), .Z(n287) );
  IVSVTX0H U564 ( .A(n287), .Z(n450) );
  ND2ASVTX2 U565 ( .A(n481), .B(n450), .Z(n475) );
  NR2ASVTX2 U566 ( .A(n481), .B(n287), .Z(n346) );
  IVSVTX2 U567 ( .A(n346), .Z(n477) );
  AO4SVTX1 U568 ( .A(n288), .B(n475), .C(n477), .D(n345), .Z(n289) );
  AO6SVTX1 U569 ( .A(n313), .B(O[27]), .C(n289), .Z(n290) );
  IVSVTX0H U570 ( .A(n309), .Z(n292) );
  AN2SVTX2 U571 ( .A(O[29]), .B(O[28]), .Z(n468) );
  AN2SVTX2 U572 ( .A(O[28]), .B(n407), .Z(n466) );
  IVSVTX0H U573 ( .A(n291), .Z(n330) );
  AO11SVTX1 U574 ( .A(n292), .B(n468), .C(n329), .D(n466), .E(n330), .F(n464), 
        .Z(n349) );
  AO11SVTX1 U575 ( .A(N[4]), .B(n321), .C(n422), .D(N[20]), .E(n423), .F(N[12]), .Z(n320) );
  AO4SVTX1 U576 ( .A(n345), .B(n475), .C(n477), .D(n320), .Z(n293) );
  AO6SVTX1 U577 ( .A(n296), .B(N[21]), .C(N[29]), .Z(n297) );
  AO7SVTX1 U578 ( .A(n394), .B(n298), .C(n297), .Z(n299) );
  AO17SVTX2 U579 ( .A(n321), .B(N[13]), .C(n299), .D(n468), .Z(n301) );
  AO3SVTX2 U580 ( .A(n302), .B(O[28]), .C(n301), .D(n300), .Z(n315) );
  IVSVTX0H U581 ( .A(n466), .Z(n453) );
  NR2ASVTX1 U582 ( .A(N[14]), .B(n319), .Z(n306) );
  AO7SVTX1 U583 ( .A(n304), .B(n404), .C(n303), .Z(n305) );
  AO1SVTX1 U584 ( .A(n307), .B(N[6]), .C(n306), .D(n305), .Z(n308) );
  AO7SVTX1 U585 ( .A(n309), .B(n453), .C(n308), .Z(n310) );
  AO6ABSVTX2 U586 ( .A(O[28]), .B(n311), .C(n310), .Z(n312) );
  AO6ABSVTX4 U587 ( .A(O[27]), .B(n315), .C(n312), .Z(n822) );
  AO2SVTX2 U588 ( .A(n313), .B(n461), .C(n346), .D(n329), .Z(n314) );
  AO7ABSVTX4 U589 ( .A(O[27]), .B(n315), .C(n314), .Z(n678) );
  IVSVTX2 U590 ( .A(n678), .Z(n768) );
  ND2SVTX2 U591 ( .A(n822), .B(n768), .Z(n819) );
  IVSVTX0H U592 ( .A(n345), .Z(n317) );
  AO11SVTX1 U593 ( .A(N[1]), .B(n321), .C(n422), .D(N[17]), .E(n423), .F(N[9]), 
        .Z(n334) );
  IVSVTX2 U594 ( .A(n334), .Z(n465) );
  AO2SVTX1 U595 ( .A(n423), .B(N[11]), .C(n422), .D(N[19]), .Z(n316) );
  AO7SVTX1 U596 ( .A(n403), .B(n319), .C(n316), .Z(n469) );
  AO11SVTX2 U597 ( .A(n317), .B(n468), .C(n465), .D(n466), .E(n469), .F(n464), 
        .Z(n325) );
  AO2SVTX1 U598 ( .A(n423), .B(N[10]), .C(n422), .D(N[18]), .Z(n318) );
  AO7SVTX1 U599 ( .A(n380), .B(n319), .C(n318), .Z(n449) );
  IVSVTX2 U600 ( .A(n320), .Z(n347) );
  AO11SVTX1 U601 ( .A(n329), .B(n468), .C(n449), .D(n466), .E(n347), .F(n464), 
        .Z(n338) );
  AO11SVTX1 U602 ( .A(N[0]), .B(n321), .C(n422), .D(N[16]), .E(n423), .F(N[8]), 
        .Z(n333) );
  AO4SVTX1 U603 ( .A(n333), .B(n475), .C(n433), .D(n477), .Z(n322) );
  AO6ABSVTX1 U604 ( .A(n481), .B(n338), .C(n322), .Z(n323) );
  AO7SVTX2 U605 ( .A(n325), .B(n284), .C(n323), .Z(n788) );
  IVSVTX2 U606 ( .A(n333), .Z(n447) );
  AO11SVTX1 U607 ( .A(n347), .B(n468), .C(n447), .D(n466), .E(n449), .F(n464), 
        .Z(n472) );
  AO2SVTX1 U608 ( .A(n423), .B(N[6]), .C(n422), .D(N[14]), .Z(n470) );
  AO4SVTX1 U609 ( .A(n477), .B(n470), .C(n433), .D(n475), .Z(n324) );
  AO7SVTX2 U610 ( .A(n472), .B(O[27]), .C(n326), .Z(n677) );
  NR2SVTX2 U611 ( .A(n788), .B(n677), .Z(n509) );
  AN2SVTX2 U612 ( .A(n422), .B(n468), .Z(n369) );
  AO2SVTX1 U613 ( .A(N[23]), .B(n369), .C(n342), .D(n468), .Z(n327) );
  AO3SVTX1 U614 ( .A(n345), .B(n435), .C(n328), .D(n327), .Z(n336) );
  AO11SVTX1 U615 ( .A(n330), .B(n468), .C(n347), .D(n466), .E(n329), .F(n464), 
        .Z(n356) );
  IVSVTX0H U616 ( .A(n475), .Z(n455) );
  AO2SVTX1 U617 ( .A(n465), .B(n346), .C(n455), .D(n449), .Z(n331) );
  AO7SVTX1 U618 ( .A(n461), .B(n356), .C(n331), .Z(n332) );
  IVSVTX0H U619 ( .A(n799), .Z(n339) );
  AO4SVTX1 U620 ( .A(n334), .B(n475), .C(n477), .D(n333), .Z(n335) );
  AO6SVTX1 U621 ( .A(n336), .B(O[27]), .C(n335), .Z(n337) );
  AO7SVTX2 U622 ( .A(O[27]), .B(n338), .C(n337), .Z(n811) );
  IVSVTX0H U623 ( .A(n811), .Z(n504) );
  AO2SVTX1 U624 ( .A(n384), .B(N[23]), .C(n342), .D(n464), .Z(n343) );
  AO3SVTX1 U625 ( .A(n345), .B(n453), .C(n344), .D(n343), .Z(n354) );
  AO2SVTX1 U626 ( .A(n347), .B(n455), .C(n346), .D(n469), .Z(n348) );
  AO7SVTX1 U627 ( .A(n461), .B(n349), .C(n348), .Z(n350) );
  IVSVTX0H U628 ( .A(n781), .Z(n357) );
  IVSVTX0H U629 ( .A(n449), .Z(n352) );
  IVSVTX0H U630 ( .A(n469), .Z(n351) );
  AO4SVTX1 U631 ( .A(n352), .B(n477), .C(n475), .D(n351), .Z(n353) );
  AO6SVTX1 U632 ( .A(O[27]), .B(n354), .C(n353), .Z(n355) );
  AO7SVTX2 U633 ( .A(n284), .B(n356), .C(n355), .Z(n786) );
  IVSVTX0H U634 ( .A(n786), .Z(n495) );
  MUX21NSVTX1 U635 ( .A(N[0]), .B(N[1]), .S(n284), .Z(n364) );
  IVSVTX0H U636 ( .A(n364), .Z(n359) );
  AN2SVTX2 U637 ( .A(n359), .B(n369), .Z(n578) );
  IVSVTX0H U638 ( .A(n578), .Z(n361) );
  NR2ASVTX1 U639 ( .A(N[0]), .B(n481), .Z(n362) );
  MUX21NSVTX1 U640 ( .A(n374), .B(n380), .S(O[27]), .Z(n370) );
  AO2SVTX1 U641 ( .A(n369), .B(n370), .C(n362), .D(n384), .Z(n572) );
  IVSVTX1 U642 ( .A(n384), .Z(n375) );
  MUX21NSVTX1 U643 ( .A(N[2]), .B(N[3]), .S(O[27]), .Z(n376) );
  NR2ASVTX2 U644 ( .A(n572), .B(n589), .Z(n365) );
  IVSVTX0H U645 ( .A(n365), .Z(n366) );
  NR2SVTX2 U646 ( .A(n367), .B(n366), .Z(n378) );
  IVSVTX0H U647 ( .A(N[4]), .Z(n379) );
  IVSVTX0H U648 ( .A(N[0]), .Z(n368) );
  AO4SVTX1 U649 ( .A(n379), .B(n381), .C(n368), .D(n405), .Z(n386) );
  IVSVTX0H U650 ( .A(n386), .Z(n373) );
  IVSVTX0H U651 ( .A(n409), .Z(n372) );
  NR2ASVTX1 U652 ( .A(N[3]), .B(O[27]), .Z(n383) );
  AO2SVTX1 U653 ( .A(n384), .B(n370), .C(n369), .D(n383), .Z(n371) );
  AO4SVTX1 U654 ( .A(n394), .B(n381), .C(n374), .D(n405), .Z(n382) );
  MUX21NSVTX1 U655 ( .A(n386), .B(n382), .S(O[27]), .Z(n391) );
  AO4SVTX2 U656 ( .A(n391), .B(n426), .C(n376), .D(n375), .Z(n599) );
  NR2SVTX1 U657 ( .A(n594), .B(n599), .Z(n377) );
  ND2SVTX2 U658 ( .A(n378), .B(n377), .Z(n568) );
  AO4SVTX1 U659 ( .A(n436), .B(n407), .C(n379), .D(n405), .Z(n395) );
  AO4SVTX1 U660 ( .A(n406), .B(n381), .C(n403), .D(n405), .Z(n390) );
  MUX21NSVTX1 U661 ( .A(n395), .B(n390), .S(n461), .Z(n399) );
  AO4SVTX1 U662 ( .A(n397), .B(n381), .C(n380), .D(n405), .Z(n389) );
  MUX21NSVTX1 U663 ( .A(n389), .B(n382), .S(n461), .Z(n388) );
  MUX21NSVTX2 U664 ( .A(n399), .B(n388), .S(n426), .Z(n609) );
  IVSVTX0H U665 ( .A(n609), .Z(n392) );
  NR2SVTX1 U666 ( .A(O[28]), .B(n481), .Z(n385) );
  AO2SVTX1 U667 ( .A(n386), .B(n385), .C(n384), .D(n383), .Z(n387) );
  AO7SVTX2 U668 ( .A(n426), .B(n388), .C(n387), .Z(n602) );
  MUX21NSVTX1 U669 ( .A(n390), .B(n389), .S(n461), .Z(n396) );
  NR2SVTX2 U670 ( .A(n602), .B(n606), .Z(n564) );
  NR2SVTX2 U671 ( .A(n568), .B(n393), .Z(n557) );
  MUX21NSVTX1 U672 ( .A(n415), .B(n395), .S(n461), .Z(n411) );
  MUX21NSVTX2 U673 ( .A(n411), .B(n396), .S(n426), .Z(n613) );
  IVSVTX0H U674 ( .A(n613), .Z(n401) );
  AO2SVTX1 U675 ( .A(n423), .B(N[2]), .C(n422), .D(N[10]), .Z(n457) );
  AO4SVTX1 U676 ( .A(n457), .B(n407), .C(n397), .D(n405), .Z(n414) );
  AO2SVTX1 U677 ( .A(n417), .B(n415), .C(n414), .D(n409), .Z(n398) );
  AO7SVTX2 U678 ( .A(O[28]), .B(n399), .C(n398), .Z(n616) );
  IVSVTX0H U679 ( .A(n616), .Z(n400) );
  IVSVTX0H U680 ( .A(N[11]), .Z(n402) );
  AO4SVTX1 U681 ( .A(n408), .B(n407), .C(n406), .D(n405), .Z(n427) );
  AO2SVTX1 U682 ( .A(n427), .B(n409), .C(n417), .D(n414), .Z(n410) );
  AO7SVTX2 U683 ( .A(O[28]), .B(n411), .C(n410), .Z(n620) );
  IVSVTX0H U684 ( .A(n620), .Z(n556) );
  AO7ABSVTX1 U685 ( .A(N[12]), .B(n422), .C(n412), .Z(n474) );
  IVSVTX0H U686 ( .A(n436), .Z(n413) );
  AO11SVTX1 U687 ( .A(n414), .B(n426), .C(n474), .D(n468), .E(n413), .F(n466), 
        .Z(n428) );
  NR2SVTX1 U688 ( .A(O[27]), .B(O[28]), .Z(n416) );
  AO2SVTX1 U689 ( .A(n427), .B(n417), .C(n416), .D(n415), .Z(n418) );
  AO7SVTX2 U690 ( .A(n461), .B(n428), .C(n418), .Z(n623) );
  IVSVTX2 U691 ( .A(n623), .Z(n419) );
  NR2SVTX2 U692 ( .A(n562), .B(n420), .Z(n421) );
  ND2SVTX2 U693 ( .A(n557), .B(n421), .Z(n527) );
  AO2SVTX1 U694 ( .A(n423), .B(N[5]), .C(n422), .D(N[13]), .Z(n476) );
  IVSVTX0H U695 ( .A(n476), .Z(n425) );
  IVSVTX0H U696 ( .A(n440), .Z(n424) );
  AO11SVTX1 U697 ( .A(n427), .B(n426), .C(n425), .D(n468), .E(n424), .F(n466), 
        .Z(n431) );
  MUX21NSVTX2 U698 ( .A(n431), .B(n428), .S(n461), .Z(n625) );
  IVSVTX0H U699 ( .A(n470), .Z(n448) );
  IVSVTX0H U700 ( .A(n457), .Z(n429) );
  AO4SVTX1 U701 ( .A(n439), .B(n461), .C(n436), .D(n475), .Z(n430) );
  AO7CSVTX2 U702 ( .A(n431), .B(O[27]), .C(n430), .Z(n628) );
  IVSVTX2 U703 ( .A(n628), .Z(n432) );
  IVSVTX0H U704 ( .A(n433), .Z(n467) );
  AO2SVTX1 U705 ( .A(n468), .B(n467), .C(n451), .D(n466), .Z(n434) );
  AO7SVTX1 U706 ( .A(n476), .B(n435), .C(n434), .Z(n442) );
  AO4SVTX1 U707 ( .A(n477), .B(n436), .C(n440), .D(n475), .Z(n437) );
  AO6SVTX1 U708 ( .A(n442), .B(O[27]), .C(n437), .Z(n438) );
  IVSVTX0H U709 ( .A(n630), .Z(n445) );
  AO11SVTX1 U710 ( .A(n447), .B(n468), .C(n474), .D(n466), .E(n448), .F(n464), 
        .Z(n458) );
  AO4SVTX1 U711 ( .A(n477), .B(n440), .C(n457), .D(n475), .Z(n441) );
  AO6SVTX1 U712 ( .A(n442), .B(n461), .C(n441), .Z(n443) );
  AO7SVTX2 U713 ( .A(n461), .B(n458), .C(n443), .Z(n637) );
  IVSVTX1 U714 ( .A(n637), .Z(n444) );
  ND2SVTX2 U715 ( .A(n445), .B(n444), .Z(n446) );
  NR2SVTX2 U716 ( .A(n546), .B(n446), .Z(n540) );
  AO11SVTX1 U717 ( .A(n449), .B(n468), .C(n448), .D(n466), .E(n447), .F(n464), 
        .Z(n483) );
  AO2SVTX1 U718 ( .A(n464), .B(n467), .C(n451), .D(n450), .Z(n452) );
  AO7SVTX1 U719 ( .A(n476), .B(n453), .C(n452), .Z(n454) );
  AO6SVTX1 U720 ( .A(n468), .B(n465), .C(n454), .Z(n460) );
  AO2ASVTX1 U721 ( .C(n455), .D(n474), .A(n460), .B(n461), .Z(n456) );
  AO7SVTX2 U722 ( .A(n461), .B(n483), .C(n456), .Z(n644) );
  AO4SVTX1 U723 ( .A(n458), .B(O[27]), .C(n457), .D(n477), .Z(n459) );
  AO7CSVTX2 U724 ( .A(n461), .B(n460), .C(n459), .Z(n641) );
  IVSVTX1 U725 ( .A(n641), .Z(n462) );
  ND2SVTX2 U726 ( .A(n463), .B(n462), .Z(n537) );
  AO11SVTX1 U727 ( .A(n469), .B(n468), .C(n467), .D(n466), .E(n465), .F(n464), 
        .Z(n480) );
  AO4SVTX1 U728 ( .A(n477), .B(n476), .C(n470), .D(n475), .Z(n471) );
  AO7SVTX2 U729 ( .A(n480), .B(O[27]), .C(n473), .Z(n651) );
  IVSVTX0H U730 ( .A(n474), .Z(n478) );
  AO4SVTX1 U731 ( .A(n478), .B(n477), .C(n476), .D(n475), .Z(n479) );
  AO7SVTX2 U732 ( .A(n483), .B(O[27]), .C(n482), .Z(n648) );
  IVSVTX1 U733 ( .A(n648), .Z(n529) );
  ND2SVTX2 U734 ( .A(n484), .B(n529), .Z(n485) );
  NR2SVTX2 U735 ( .A(n537), .B(n485), .Z(n486) );
  ND2SVTX2 U736 ( .A(n540), .B(n486), .Z(n487) );
  NR2SVTX2 U737 ( .A(n527), .B(n487), .Z(n523) );
  IVSVTX4 U738 ( .A(n523), .Z(n533) );
  NR2SVTX2 U739 ( .A(n488), .B(n533), .Z(n491) );
  ND2SVTX2 U740 ( .A(n822), .B(n678), .Z(n782) );
  IVSVTX2 U741 ( .A(n782), .Z(n494) );
  IVSVTX2 U742 ( .A(n214), .Z(n793) );
  NR2SVTX2 U743 ( .A(n781), .B(n779), .Z(n812) );
  IVSVTX2 U744 ( .A(n507), .Z(n500) );
  ND2SVTX2 U745 ( .A(n495), .B(n500), .Z(n496) );
  NR2SVTX2 U746 ( .A(n496), .B(n533), .Z(n497) );
  ENSVTX1 U747 ( .A(n781), .B(n497), .Z(n515) );
  BFSVTX2 U748 ( .A(n498), .Z(n656) );
  IVSVTX0H U749 ( .A(n499), .Z(n501) );
  ND2SVTX2 U750 ( .A(n501), .B(n500), .Z(n502) );
  NR2SVTX2 U751 ( .A(n502), .B(n533), .Z(n503) );
  ENSVTX1 U752 ( .A(n773), .B(n503), .Z(n657) );
  AO11NSVTX2 U753 ( .A(n781), .B(n659), .C(n658), .D(n515), .E(n656), .F(n657), 
        .Z(n798) );
  NR2SVTX2 U754 ( .A(n505), .B(n533), .Z(n506) );
  ENSVTX1 U755 ( .A(n799), .B(n506), .Z(n512) );
  NR2SVTX2 U756 ( .A(n507), .B(n533), .Z(n508) );
  ENSVTX1 U757 ( .A(n786), .B(n508), .Z(n516) );
  AO11NSVTX2 U758 ( .A(n799), .B(n659), .C(n658), .D(n512), .E(n656), .F(n516), 
        .Z(n787) );
  NR2SVTX2 U759 ( .A(n788), .B(n787), .Z(n522) );
  IVSVTX0H U760 ( .A(n509), .Z(n510) );
  NR2SVTX2 U761 ( .A(n510), .B(n533), .Z(n511) );
  AO11NSVTX2 U762 ( .A(n811), .B(n659), .C(n658), .D(n526), .E(n656), .F(n512), 
        .Z(n676) );
  ND2SVTX2 U763 ( .A(n677), .B(n676), .Z(n514) );
  ND2SVTX2 U764 ( .A(n788), .B(n787), .Z(n513) );
  AO11NSVTX2 U765 ( .A(n786), .B(n659), .C(n658), .D(n516), .E(n656), .F(n515), 
        .Z(n810) );
  NR2SVTX2 U766 ( .A(n811), .B(n810), .Z(n521) );
  IVSVTX1 U767 ( .A(n521), .Z(n518) );
  ND2SVTX2 U768 ( .A(n799), .B(n798), .Z(n666) );
  AO7SVTX1 U769 ( .A(n664), .B(n667), .C(n666), .Z(n654) );
  NR2SVTX2 U770 ( .A(n677), .B(n676), .Z(n520) );
  NR3SVTX2 U771 ( .A(n522), .B(n521), .C(n520), .Z(n668) );
  IVSVTX1 U772 ( .A(n668), .Z(n652) );
  IVSVTX0H U773 ( .A(n677), .Z(n524) );
  ND2SVTX2 U774 ( .A(n524), .B(n523), .Z(n525) );
  EOSVTX1 U775 ( .A(n788), .B(n525), .Z(n645) );
  IVSVTX4 U776 ( .A(n527), .Z(n560) );
  IVSVTX0H U777 ( .A(n537), .Z(n528) );
  IVSVTX0H U778 ( .A(n540), .Z(n536) );
  NR2SVTX1 U779 ( .A(n530), .B(n536), .Z(n531) );
  ND2SVTX2 U780 ( .A(n560), .B(n531), .Z(n532) );
  EOSVTX1 U781 ( .A(n651), .B(n532), .Z(n638) );
  EOSVTX1 U782 ( .A(n677), .B(n533), .Z(n646) );
  NR2SVTX1 U783 ( .A(n641), .B(n536), .Z(n534) );
  ND2SVTX2 U784 ( .A(n560), .B(n534), .Z(n535) );
  EOSVTX2 U785 ( .A(n644), .B(n535), .Z(n542) );
  NR2SVTX1 U786 ( .A(n537), .B(n536), .Z(n538) );
  ND2SVTX2 U787 ( .A(n560), .B(n538), .Z(n539) );
  EOSVTX1 U788 ( .A(n648), .B(n539), .Z(n639) );
  NR2SVTX2 U789 ( .A(n637), .B(n636), .Z(n697) );
  ND2SVTX2 U790 ( .A(n540), .B(n560), .Z(n541) );
  AO11NSVTX4 U791 ( .A(n641), .B(n659), .C(n658), .D(n545), .E(n656), .F(n542), 
        .Z(n629) );
  NR2SVTX2 U792 ( .A(n630), .B(n629), .Z(n632) );
  IVSVTX2 U793 ( .A(n632), .Z(n711) );
  NR2SVTX2 U794 ( .A(n630), .B(n546), .Z(n543) );
  ND2SVTX2 U795 ( .A(n543), .B(n560), .Z(n544) );
  AO11NSVTX2 U796 ( .A(n637), .B(n793), .C(n494), .D(n549), .E(n656), .F(n545), 
        .Z(n627) );
  NR2SVTX2 U797 ( .A(n628), .B(n627), .Z(n702) );
  IVSVTX0H U798 ( .A(n546), .Z(n547) );
  ND2SVTX2 U799 ( .A(n547), .B(n560), .Z(n548) );
  AO11NSVTX2 U800 ( .A(n630), .B(n793), .C(n658), .D(n552), .E(n656), .F(n549), 
        .Z(n624) );
  NR2SVTX2 U801 ( .A(n625), .B(n624), .Z(n705) );
  ND2SVTX2 U802 ( .A(n550), .B(n560), .Z(n551) );
  AO11NSVTX2 U803 ( .A(n628), .B(n793), .C(n494), .D(n618), .E(n656), .F(n552), 
        .Z(n622) );
  ND3ABSVTX2 U804 ( .A(n702), .B(n705), .C(n718), .Z(n713) );
  IVSVTX0H U805 ( .A(n713), .Z(n554) );
  AN2SVTX2 U806 ( .A(n711), .B(n554), .Z(n634) );
  IVSVTX0H U807 ( .A(n562), .Z(n555) );
  IVSVTX2 U808 ( .A(n557), .Z(n566) );
  NR2SVTX2 U809 ( .A(n558), .B(n566), .Z(n559) );
  ENSVTX1 U810 ( .A(n623), .B(n559), .Z(n610) );
  ENSVTX1 U811 ( .A(n625), .B(n560), .Z(n617) );
  ENSVTX1 U812 ( .A(n616), .B(n561), .Z(n603) );
  NR2SVTX2 U813 ( .A(n562), .B(n566), .Z(n563) );
  ENSVTX1 U814 ( .A(n620), .B(n563), .Z(n611) );
  NR2SVTX2 U815 ( .A(n609), .B(n608), .Z(n736) );
  NR2ASVTX1 U816 ( .A(n564), .B(n568), .Z(n565) );
  ENSVTX1 U817 ( .A(n609), .B(n565), .Z(n595) );
  EOSVTX1 U818 ( .A(n613), .B(n566), .Z(n604) );
  NR2SVTX2 U819 ( .A(n602), .B(n601), .Z(n744) );
  IVSVTX0H U820 ( .A(n568), .Z(n567) );
  IVSVTX0H U821 ( .A(n606), .Z(n571) );
  IVSVTX0H U822 ( .A(n602), .Z(n569) );
  NR2ASVTX1 U823 ( .A(n569), .B(n568), .Z(n570) );
  EOSVTX1 U824 ( .A(n571), .B(n570), .Z(n597) );
  AO11NSVTX2 U825 ( .A(n602), .B(n793), .C(n658), .D(n586), .E(n498), .F(n597), 
        .Z(n593) );
  NR2SVTX2 U826 ( .A(n594), .B(n593), .Z(n753) );
  IVSVTX0H U827 ( .A(n572), .Z(n582) );
  IVSVTX0H U828 ( .A(n594), .Z(n573) );
  IVSVTX0H U829 ( .A(n599), .Z(n587) );
  AO11NSVTX1 U830 ( .A(n594), .B(n793), .C(n494), .D(n573), .E(n498), .F(n587), 
        .Z(n581) );
  NR2SVTX2 U831 ( .A(n582), .B(n581), .Z(n585) );
  IVSVTX0H U832 ( .A(n589), .Z(n574) );
  AO11NSVTX2 U833 ( .A(n589), .B(n793), .C(n494), .D(n574), .E(n498), .F(n573), 
        .Z(n577) );
  AN2SVTX2 U834 ( .A(n578), .B(n577), .Z(n579) );
  ND2SVTX2 U835 ( .A(n582), .B(n581), .Z(n583) );
  AO11NSVTX4 U836 ( .A(n599), .B(n793), .C(n658), .D(n587), .E(n498), .F(n586), 
        .Z(n588) );
  OR2SVTX2 U837 ( .A(n589), .B(n588), .Z(n591) );
  AN2SVTX2 U838 ( .A(n589), .B(n588), .Z(n590) );
  ND2SVTX2 U839 ( .A(n594), .B(n593), .Z(n755) );
  AO2SVTX1 U840 ( .A(n595), .B(n498), .C(n606), .D(n793), .Z(n596) );
  OR2SVTX2 U841 ( .A(n599), .B(n598), .Z(n749) );
  ND2SVTX2 U842 ( .A(n599), .B(n598), .Z(n750) );
  IVSVTX0H U843 ( .A(n750), .Z(n600) );
  ND2SVTX2 U844 ( .A(n602), .B(n601), .Z(n746) );
  AO11NSVTX2 U845 ( .A(n613), .B(n793), .C(n658), .D(n604), .E(n656), .F(n603), 
        .Z(n605) );
  ND2SVTX2 U846 ( .A(n606), .B(n605), .Z(n741) );
  IVSVTX0H U847 ( .A(n741), .Z(n607) );
  AO11NSVTX2 U848 ( .A(n620), .B(n793), .C(n494), .D(n611), .E(n656), .F(n610), 
        .Z(n612) );
  OR2SVTX2 U849 ( .A(n613), .B(n612), .Z(n732) );
  ND2SVTX2 U850 ( .A(n613), .B(n612), .Z(n733) );
  IVSVTX0H U851 ( .A(n733), .Z(n614) );
  IVSVTX0H U852 ( .A(n724), .Z(n621) );
  AO6SVTX8 U853 ( .A(n725), .B(n723), .C(n621), .Z(n720) );
  ND2SVTX2 U854 ( .A(n623), .B(n622), .Z(n719) );
  ND2SVTX2 U855 ( .A(n625), .B(n624), .Z(n717) );
  IVSVTX0H U856 ( .A(n717), .Z(n626) );
  AO6ABSVTX2 U857 ( .A(n705), .B(n719), .C(n626), .Z(n707) );
  ND2SVTX1 U858 ( .A(n628), .B(n627), .Z(n704) );
  ND2SVTX2 U859 ( .A(n630), .B(n629), .Z(n712) );
  IVSVTX0H U860 ( .A(n712), .Z(n631) );
  AO7ASVTX8 U861 ( .A(n634), .B(n720), .C(n633), .Z(n635) );
  IVSVTX6 U862 ( .A(n635), .Z(n700) );
  ND2SVTX2 U863 ( .A(n637), .B(n636), .Z(n699) );
  AO7SVTX8 U864 ( .A(n697), .B(n700), .C(n699), .Z(n845) );
  AO11NSVTX4 U865 ( .A(n648), .B(n659), .C(n658), .D(n639), .E(n656), .F(n638), 
        .Z(n640) );
  OR2SVTX2 U866 ( .A(n641), .B(n640), .Z(n843) );
  ND2SVTX1 U867 ( .A(n641), .B(n640), .Z(n844) );
  AO6SVTX8 U868 ( .A(n845), .B(n843), .C(n642), .Z(n766) );
  ND2SVTX1 U869 ( .A(n644), .B(n643), .Z(n765) );
  AO7SVTX8 U870 ( .A(n763), .B(n766), .C(n765), .Z(n695) );
  AO11NSVTX2 U871 ( .A(n677), .B(n659), .C(n658), .D(n646), .E(n656), .F(n645), 
        .Z(n647) );
  OR2SVTX2 U872 ( .A(n648), .B(n647), .Z(n693) );
  ND2SVTX2 U873 ( .A(n648), .B(n647), .Z(n694) );
  IVSVTX0H U874 ( .A(n694), .Z(n649) );
  AO6SVTX8 U875 ( .A(n695), .B(n693), .C(n649), .Z(n761) );
  ND2SVTX2 U876 ( .A(n786), .B(n785), .Z(n681) );
  AO6SVTX8 U877 ( .A(n682), .B(n680), .C(n660), .Z(n815) );
  ND2SVTX2 U878 ( .A(n781), .B(n779), .Z(n814) );
  ND2ASVTX8 U879 ( .A(n789), .B(n794), .Z(n817) );
  IVSVTX0H U880 ( .A(n822), .Z(n679) );
  ND3SVTX1 U881 ( .A(n794), .B(n817), .C(n679), .Z(n663) );
  OR2SVTX2 U882 ( .A(n673), .B(n672), .Z(n689) );
  IVSVTX0H U883 ( .A(n664), .Z(n665) );
  EOSVTX1 U884 ( .A(n670), .B(n669), .Z(n671) );
  ND2SVTX2 U885 ( .A(n673), .B(n672), .Z(n690) );
  ND2ASVTX2 U886 ( .A(n822), .B(n678), .Z(n805) );
  AO7SVTX1 U887 ( .A(n789), .B(n679), .C(n805), .Z(n827) );
  ENSVTX1 U888 ( .A(n683), .B(n682), .Z(n684) );
  NR2ASVTX2 U889 ( .A(n684), .B(n817), .Z(n826) );
  ND2SVTX2 U890 ( .A(n686), .B(n685), .Z(n832) );
  NR2SVTX2 U891 ( .A(n686), .B(n685), .Z(n834) );
  IVSVTX0H U892 ( .A(n834), .Z(n687) );
  EOSVTX1 U893 ( .A(n833), .B(n688), .Z(O[18]) );
  ENSVTX1 U894 ( .A(n692), .B(n691), .Z(O[17]) );
  ENSVTX1 U895 ( .A(n696), .B(n695), .Z(O[15]) );
  IVSVTX0H U896 ( .A(n697), .Z(n698) );
  EOSVTX1 U897 ( .A(n701), .B(n700), .Z(O[12]) );
  IVSVTX0H U898 ( .A(n702), .Z(n703) );
  IVSVTX0H U899 ( .A(n705), .Z(n716) );
  NR2ASVTX1 U900 ( .A(n707), .B(n706), .Z(n708) );
  EOSVTX1 U901 ( .A(n709), .B(n708), .Z(O[10]) );
  EOSVTX1 U902 ( .A(n710), .B(n720), .Z(O[8]) );
  ND2SVTX1 U903 ( .A(n712), .B(n711), .Z(n715) );
  AO7SVTX1 U904 ( .A(n713), .B(n720), .C(n212), .Z(n714) );
  ENSVTX1 U905 ( .A(n715), .B(n714), .Z(O[11]) );
  AO7SVTX1 U906 ( .A(n553), .B(n720), .C(n719), .Z(n721) );
  ENSVTX1 U907 ( .A(n722), .B(n721), .Z(O[9]) );
  ENSVTX1 U908 ( .A(n726), .B(n725), .Z(O[7]) );
  IVSVTX0H U909 ( .A(n727), .Z(n728) );
  EOSVTX1 U910 ( .A(n731), .B(n730), .Z(O[6]) );
  ENSVTX1 U911 ( .A(n735), .B(n734), .Z(O[5]) );
  IVSVTX0H U912 ( .A(n736), .Z(n737) );
  EOSVTX1 U913 ( .A(n740), .B(n739), .Z(O[4]) );
  ND2SVTX1 U914 ( .A(n741), .B(n211), .Z(n743) );
  ENSVTX1 U915 ( .A(n743), .B(n742), .Z(O[3]) );
  IVSVTX0H U916 ( .A(n744), .Z(n745) );
  ND2SVTX1 U917 ( .A(n746), .B(n745), .Z(n748) );
  EOSVTX1 U918 ( .A(n748), .B(n747), .Z(O[2]) );
  ND2SVTX1 U919 ( .A(n750), .B(n749), .Z(n752) );
  ENSVTX1 U920 ( .A(n752), .B(n751), .Z(O[1]) );
  IVSVTX0H U921 ( .A(n753), .Z(n754) );
  ND2SVTX1 U922 ( .A(n755), .B(n754), .Z(n757) );
  EOSVTX1 U923 ( .A(n757), .B(n756), .Z(O[0]) );
  IVSVTX0H U924 ( .A(n758), .Z(n759) );
  EOSVTX1 U925 ( .A(n762), .B(n761), .Z(O[16]) );
  IVSVTX0H U926 ( .A(n763), .Z(n764) );
  EOSVTX1 U927 ( .A(n767), .B(n766), .Z(O[14]) );
  AO7SVTX1 U928 ( .A(n782), .B(n775), .C(n214), .Z(n769) );
  AO6SVTX1 U929 ( .A(n789), .B(n768), .C(n662), .Z(n804) );
  EOSVTX1 U930 ( .A(n769), .B(n770), .Z(n836) );
  IVSVTX2 U931 ( .A(n817), .Z(n821) );
  FA1SVTX1 U932 ( .A(n773), .B(n772), .CI(n771), .CO(n777), .Z(n784) );
  FA1SVTX1 U933 ( .A(n778), .B(n777), .CI(n776), .CO(n851), .Z(n848) );
  FA1SVTX1 U934 ( .A(n781), .B(n780), .CI(n779), .CO(n771), .Z(n796) );
  NR2ASVTX1 U935 ( .A(n782), .B(n817), .Z(n795) );
  HA1SVTX1 U936 ( .A(n786), .B(n785), .CO(n780), .S(n808) );
  HA1SVTX1 U937 ( .A(n788), .B(n787), .CO(n809), .S(n828) );
  IVSVTX0H U938 ( .A(n805), .Z(n790) );
  AO7SVTX1 U939 ( .A(n790), .B(n498), .C(n789), .Z(n791) );
  AO3SVTX1 U940 ( .A(n794), .B(n793), .C(n792), .D(n791), .Z(n806) );
  FA1SVTX1 U941 ( .A(n796), .B(n821), .CI(n795), .CO(n857), .Z(n853) );
  FA1SVTX1 U942 ( .A(n799), .B(n798), .CI(n797), .CO(n807), .Z(n825) );
  IVSVTX0H U943 ( .A(n800), .Z(n802) );
  ENSVTX1 U944 ( .A(n802), .B(n801), .Z(n803) );
  NR2ASVTX1 U945 ( .A(n803), .B(n817), .Z(n824) );
  AO3SVTX1 U946 ( .A(n817), .B(n805), .C(n804), .D(n819), .Z(n823) );
  FA1SVTX1 U947 ( .A(n808), .B(n807), .CI(n806), .CO(n854), .Z(n859) );
  FA1SVTX1 U948 ( .A(n811), .B(n810), .CI(n809), .CO(n797), .Z(n831) );
  IVSVTX0H U949 ( .A(n812), .Z(n813) );
  NR2ASVTX1 U950 ( .A(n818), .B(n817), .Z(n830) );
  FA1SVTX1 U951 ( .A(n825), .B(n824), .CI(n823), .CO(n860), .Z(n841) );
  EOSVTX4 U952 ( .A(n836), .B(n835), .Z(O[26]) );
  FA1SVTX4 U953 ( .A(n842), .B(n841), .CI(n840), .CO(n858), .Z(O[20]) );
  ND2SVTX1 U954 ( .A(n844), .B(n843), .Z(n846) );
  ENSVTX1 U955 ( .A(n846), .B(n845), .Z(O[13]) );
endmodule

