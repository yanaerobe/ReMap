
module m_rangemapping ( N, O );
  input [31:0] N;
  output [31:0] O;
  wire   n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917;

  ENSVTX1 U296 ( .A(n808), .B(n807), .Z(O[24]) );
  EOSVTX1 U297 ( .A(n827), .B(n826), .Z(O[21]) );
  ENSVTX0H U298 ( .A(n910), .B(n909), .Z(O[20]) );
  EOSVTX0H U299 ( .A(n822), .B(n821), .Z(O[19]) );
  ENSVTX0H U300 ( .A(n817), .B(n816), .Z(O[22]) );
  IVSVTX0H U301 ( .A(n214), .Z(n804) );
  IVSVTX0H U302 ( .A(n869), .Z(n886) );
  F_FA1SVTX1 U303 ( .A(n799), .B(n798), .CI(n797), .CO(n700), .Z(n805) );
  IVSVTX0H U304 ( .A(n707), .Z(n798) );
  OR2SVTX2 U305 ( .A(n793), .B(n792), .Z(n814) );
  F_FA1SVTX1 U306 ( .A(n706), .B(n705), .CI(n704), .CO(n797), .Z(n802) );
  AO7SVTX4 U307 ( .A(n822), .B(n818), .C(n820), .Z(n909) );
  NR2ASVTX1 U308 ( .A(n912), .B(n771), .Z(n790) );
  AO7SVTX1 U309 ( .A(n742), .B(n719), .C(n718), .Z(n787) );
  NR2ASVTX1 U310 ( .A(n772), .B(n771), .Z(n775) );
  NR2ASVTX1 U311 ( .A(n741), .B(n771), .Z(n745) );
  IVSVTX0H U312 ( .A(n731), .Z(n709) );
  F_FA1SVTX1 U313 ( .A(n757), .B(n756), .CI(n755), .CO(n721), .Z(n777) );
  EOSVTX0H U314 ( .A(n740), .B(n767), .Z(n741) );
  IVSVTX0H U315 ( .A(n697), .Z(n742) );
  IVSVTX0H U316 ( .A(n760), .Z(n744) );
  NR2SVTX2 U317 ( .A(n618), .B(n696), .Z(n697) );
  AO2NSVTX1 U318 ( .A(n672), .B(n661), .C(n650), .D(n717), .Z(n704) );
  IVSVTX0H U319 ( .A(n649), .Z(n650) );
  EOSVTX1 U320 ( .A(n648), .B(n649), .Z(n661) );
  EOSVTX1 U321 ( .A(n799), .B(n653), .Z(n660) );
  EOSVTX0H U322 ( .A(n706), .B(n655), .Z(n659) );
  EOSVTX1 U323 ( .A(n715), .B(n666), .Z(n686) );
  EOSVTX0H U324 ( .A(n737), .B(n439), .Z(n444) );
  AO3SVTX1 U325 ( .A(n623), .B(n640), .C(n600), .D(n599), .Z(n799) );
  F_MUX21NSVTX0H U326 ( .A(n603), .B(n598), .S(O[27]), .Z(n600) );
  IVSVTX0H U327 ( .A(n877), .Z(n884) );
  AO7SVTX2 U328 ( .A(n903), .B(n907), .C(n905), .Z(n895) );
  EOSVTX1 U329 ( .A(n559), .B(n530), .Z(n557) );
  AO11NSVTX1 U330 ( .A(n672), .B(n490), .C(n689), .D(n508), .E(n497), .F(n717), 
        .Z(n498) );
  F_MUX21NSVTX0H U331 ( .A(n603), .B(n612), .S(n274), .Z(n605) );
  IVSVTX2 U332 ( .A(n911), .Z(n689) );
  MUX21NSVTX1 U333 ( .A(n575), .B(n320), .S(n274), .Z(n322) );
  IVSVTX2 U334 ( .A(n911), .Z(n719) );
  IVSVTX0H U335 ( .A(n641), .Z(n266) );
  ND2SVTX2 U336 ( .A(n760), .B(n648), .Z(n912) );
  IVSVTX0H U337 ( .A(n429), .Z(n415) );
  IVSVTX0H U338 ( .A(n423), .Z(n394) );
  F_MUX21NSVTX1 U339 ( .A(N[0]), .B(N[1]), .S(O[27]), .Z(n349) );
  F_MUX21NSVTX1 U340 ( .A(n368), .B(n362), .S(n274), .Z(n379) );
  IVSVTX2 U341 ( .A(n630), .Z(n640) );
  AN2BSVTX2 U342 ( .A(n344), .B(n374), .Z(n377) );
  F_ND2ASVTX2 U343 ( .A(O[27]), .B(n326), .Z(n633) );
  IVSVTX6 U344 ( .A(O[27]), .Z(n274) );
  AO2SVTX1 U345 ( .A(n421), .B(n288), .C(n571), .D(n595), .Z(n289) );
  AO1SVTX1 U346 ( .A(n366), .B(n601), .C(n300), .D(n299), .Z(n316) );
  NR2ASVTX2 U347 ( .A(n366), .B(O[28]), .Z(n326) );
  IVSVTX2 U348 ( .A(n622), .Z(n421) );
  AO21SVTX1 U349 ( .A(N[22]), .B(n271), .C(n260), .D(n221), .Z(n241) );
  ND2ASVTX4 U350 ( .A(O[29]), .B(O[28]), .Z(n626) );
  AO21SVTX1 U351 ( .A(N[6]), .B(n365), .C(n262), .D(n226), .Z(n229) );
  IVSVTX0H U352 ( .A(N[21]), .Z(n271) );
  AO7SVTX1 U353 ( .A(n313), .B(n260), .C(n250), .Z(n259) );
  AO6SVTX1 U354 ( .A(n245), .B(n244), .C(n243), .Z(n249) );
  IVSVTX0H U355 ( .A(N[22]), .Z(n313) );
  IVSVTX0H U356 ( .A(N[16]), .Z(n227) );
  IVSVTX2 U357 ( .A(N[14]), .Z(n315) );
  IVSVTX0H U358 ( .A(n561), .Z(n418) );
  F_ND2SVTX0H U359 ( .A(N[0]), .B(n306), .Z(n292) );
  ND3SVTX1 U360 ( .A(n274), .B(N[3]), .C(n572), .Z(n341) );
  B_ND2SVTX0H U361 ( .A(n762), .B(n761), .Z(n770) );
  AO6ASVTX1 U362 ( .A(n361), .B(n306), .C(n304), .Z(n602) );
  AO11NSVTX2 U363 ( .A(n715), .B(n689), .C(n445), .D(n688), .E(n687), .F(n686), 
        .Z(n755) );
  EOSVTX2 U364 ( .A(n521), .B(n461), .Z(n506) );
  EOSVTX1 U365 ( .A(n551), .B(n452), .Z(n542) );
  EOSVTX2 U366 ( .A(n757), .B(n580), .Z(n673) );
  AO3SVTX1 U367 ( .A(n625), .B(n633), .C(n605), .D(n604), .Z(n706) );
  AO11NSVTX1 U368 ( .A(n501), .B(n719), .C(n717), .D(n490), .E(n672), .F(n466), 
        .Z(n487) );
  OR2SVTX1 U369 ( .A(n431), .B(n430), .Z(n551) );
  IVSVTX0H U370 ( .A(N[1]), .Z(n347) );
  IVSVTX0H U371 ( .A(n231), .Z(n251) );
  EOSVTX0H U372 ( .A(n874), .B(n873), .Z(O[8]) );
  ENSVTX0H U373 ( .A(n831), .B(n830), .Z(O[18]) );
  B_ND2SVTX1 U374 ( .A(n806), .B(n805), .Z(n808) );
  B_ND2SVTX1 U375 ( .A(n834), .B(n833), .Z(n835) );
  B_ND2SVTX2 U376 ( .A(n785), .B(n784), .Z(n825) );
  NR2SVTX2 U377 ( .A(n785), .B(n784), .Z(n823) );
  ND2SVTX6 U378 ( .A(n710), .B(n711), .Z(n696) );
  B_ND2SVTX0H U379 ( .A(n723), .B(n764), .Z(n725) );
  B_ND2SVTX2 U380 ( .A(n669), .B(n647), .Z(n649) );
  B_ND2SVTX2 U381 ( .A(n540), .B(n451), .Z(n452) );
  B_ND2SVTX2 U382 ( .A(n669), .B(n665), .Z(n666) );
  B_ND2SVTX2 U383 ( .A(n670), .B(n669), .Z(n671) );
  BFSVTX6 U384 ( .A(n687), .Z(n672) );
  F_ND2SVTX1 U385 ( .A(n642), .B(n663), .Z(n643) );
  MUX21NSVTX2 U386 ( .A(n317), .B(n598), .S(n274), .Z(n318) );
  CTIVSVTX2 U387 ( .A(n521), .Z(n390) );
  IVSVTX2 U388 ( .A(n510), .Z(n493) );
  B_ND2SVTX1 U389 ( .A(n421), .B(n637), .Z(n327) );
  IVSVTX4 U390 ( .A(n626), .Z(n571) );
  NR3ABSVTX6 U391 ( .A(n238), .B(n237), .C(n236), .Z(n389) );
  B_IVSVTX1 U392 ( .A(N[9]), .Z(n286) );
  CTIVSVTX2 U393 ( .A(N[5]), .Z(n365) );
  B_ND2SVTX2 U394 ( .A(n825), .B(n824), .Z(n827) );
  AO6SVTX4 U395 ( .A(n828), .B(n831), .C(n751), .Z(n822) );
  B_ND2SVTX2 U396 ( .A(n908), .B(n213), .Z(n910) );
  B_ND2SVTX2 U397 ( .A(n793), .B(n792), .Z(n815) );
  B_ND2SVTX2 U398 ( .A(n774), .B(n773), .Z(n820) );
  ND3SVTX2 U399 ( .A(n742), .B(n771), .C(n744), .Z(n743) );
  F_ND2ASVTX2 U400 ( .A(n716), .B(n708), .Z(n913) );
  AO7CSVTX2 U401 ( .A(n789), .B(n760), .C(n759), .Z(n776) );
  B_ND2SVTX2 U402 ( .A(n709), .B(n789), .Z(n707) );
  IVSVTX4 U403 ( .A(n789), .Z(n771) );
  AO6SVTX2 U404 ( .A(n698), .B(n729), .C(n697), .Z(n708) );
  IVSVTX2 U405 ( .A(n729), .Z(n211) );
  F_ND2ASVTX1 U406 ( .A(n733), .B(n732), .Z(n736) );
  AO7SVTX2 U407 ( .A(n870), .B(n526), .C(n525), .Z(n527) );
  B_ND2SVTX2 U408 ( .A(n847), .B(n850), .Z(n556) );
  AO6SVTX4 U409 ( .A(n895), .B(n503), .C(n502), .Z(n591) );
  B_ND2SVTX1 U410 ( .A(n839), .B(n838), .Z(n846) );
  IVSVTX2 U411 ( .A(n693), .Z(n764) );
  AO7SVTX2 U412 ( .A(n678), .B(n585), .C(n677), .Z(n733) );
  B_ND2SVTX1 U413 ( .A(n859), .B(n858), .Z(n861) );
  B_ND2SVTX2 U414 ( .A(n546), .B(n545), .Z(n859) );
  AO6SVTX2 U415 ( .A(n486), .B(n485), .C(n484), .Z(n907) );
  OR2SVTX4 U416 ( .A(n706), .B(n704), .Z(n710) );
  B_ND2SVTX1 U417 ( .A(n881), .B(n880), .Z(n883) );
  B_ND2SVTX1 U418 ( .A(n590), .B(n589), .Z(n594) );
  B_ND2SVTX2 U419 ( .A(n529), .B(n669), .Z(n530) );
  F_ND2SVTX1 U420 ( .A(n669), .B(n654), .Z(n655) );
  B_ND2SVTX1 U421 ( .A(n889), .B(n888), .Z(n891) );
  B_ND2SVTX2 U422 ( .A(n442), .B(n669), .Z(n443) );
  F_ENSVTX2 U423 ( .A(n564), .B(n669), .Z(n536) );
  B_ND2SVTX2 U424 ( .A(n669), .B(n652), .Z(n653) );
  B_ND2SVTX1 U425 ( .A(n478), .B(n477), .Z(n479) );
  B_ND2SVTX2 U426 ( .A(n450), .B(n540), .Z(n446) );
  F_ND2SVTX1 U427 ( .A(n672), .B(n462), .Z(n458) );
  B_ND2SVTX2 U428 ( .A(n645), .B(n644), .Z(n656) );
  BFSVTX8 U429 ( .A(n445), .Z(n717) );
  F_ND2SVTX1 U430 ( .A(n618), .B(n617), .Z(n646) );
  B_ND2SVTX2 U431 ( .A(n456), .B(n540), .Z(n457) );
  F_ND2SVTX1 U432 ( .A(n663), .B(n662), .Z(n664) );
  IVSVTX4 U433 ( .A(n912), .Z(n687) );
  IVSVTX4 U434 ( .A(n447), .Z(n540) );
  B_ND2SVTX2 U435 ( .A(n529), .B(n331), .Z(n441) );
  AO7SVTX4 U436 ( .A(n401), .B(n400), .C(n399), .Z(n523) );
  B_ND2SVTX2 U437 ( .A(n433), .B(n432), .Z(n538) );
  F_ND2SVTX1 U438 ( .A(n493), .B(n492), .Z(n494) );
  IVSVTX2 U439 ( .A(n799), .Z(n618) );
  MUX21NSVTX2 U440 ( .A(n398), .B(n397), .S(n274), .Z(n399) );
  CTIVSVTX2 U441 ( .A(n757), .Z(n619) );
  CTIVSVTX2 U442 ( .A(n559), .Z(n331) );
  ND2ASVTX4 U443 ( .A(n319), .B(n318), .Z(n648) );
  CTIVSVTX2 U444 ( .A(n722), .Z(n663) );
  IVSVTX2 U445 ( .A(n464), .Z(n495) );
  MUX21NSVTX1 U446 ( .A(n628), .B(n634), .S(n274), .Z(n632) );
  MUX21NSVTX1 U447 ( .A(n628), .B(n612), .S(O[27]), .Z(n614) );
  CTIVSVTX2 U448 ( .A(n551), .Z(n432) );
  IVSVTX2 U449 ( .A(n317), .Z(n311) );
  MUX21NSVTX1 U450 ( .A(n334), .B(n333), .S(O[27]), .Z(n336) );
  B_ND2SVTX2 U451 ( .A(n463), .B(n212), .Z(n356) );
  AO7SVTX2 U452 ( .A(n596), .B(n379), .C(n378), .Z(n501) );
  MUX21NSVTX2 U453 ( .A(n385), .B(n379), .S(n596), .Z(n510) );
  MUX21NSVTX1 U454 ( .A(n333), .B(n320), .S(O[27]), .Z(n272) );
  B_ND2SVTX1 U455 ( .A(n413), .B(n636), .Z(n321) );
  B_ND2SVTX1 U456 ( .A(n420), .B(n630), .Z(n416) );
  NR2SVTX2 U457 ( .A(n349), .B(n351), .Z(n473) );
  MUX21NSVTX1 U458 ( .A(n377), .B(n376), .S(O[27]), .Z(n378) );
  F_ND2SVTX1 U459 ( .A(n606), .B(n636), .Z(n599) );
  B_ND2SVTX1 U460 ( .A(n422), .B(n630), .Z(n335) );
  AO4SVTX2 U461 ( .A(n364), .B(n340), .C(n357), .D(n359), .Z(n375) );
  IVSVTX4 U462 ( .A(n624), .Z(n570) );
  AO2SVTX2 U463 ( .A(n384), .B(N[10]), .C(n363), .D(N[2]), .Z(n409) );
  F_MUX21NSVTX1 U464 ( .A(N[1]), .B(N[2]), .S(O[27]), .Z(n350) );
  B_ND2SVTX2 U465 ( .A(N[23]), .B(n387), .Z(n280) );
  IVSVTX4 U466 ( .A(O[28]), .Z(n596) );
  ND2ASVTX6 U467 ( .A(n366), .B(O[28]), .Z(n622) );
  OR2SVTX6 U468 ( .A(n366), .B(O[28]), .Z(n624) );
  B_ND2SVTX1 U469 ( .A(N[5]), .B(n306), .Z(n283) );
  CTIVSVTX2 U470 ( .A(n306), .Z(n298) );
  NR2SVTX2 U471 ( .A(O[31]), .B(n263), .Z(n306) );
  AO7ASVTX6 U472 ( .A(n262), .B(O[31]), .C(n261), .Z(n263) );
  B_ND2SVTX2 U473 ( .A(N[19]), .B(n231), .Z(n238) );
  AO1SVTX2 U474 ( .A(n359), .B(N[27]), .C(N[31]), .D(n232), .Z(n237) );
  ND2SVTX6 U475 ( .A(n217), .B(n359), .Z(n260) );
  NR2SVTX1 U476 ( .A(N[30]), .B(n218), .Z(n219) );
  CTIVSVTX2 U477 ( .A(N[6]), .Z(n360) );
  NR2ASVTX4 U478 ( .A(n214), .B(n915), .Z(n916) );
  AO6SVTX6 U479 ( .A(n807), .B(n805), .C(n803), .Z(n915) );
  AO7SVTX6 U480 ( .A(n809), .B(n812), .C(n811), .Z(n807) );
  AO6SVTX6 U481 ( .A(n816), .B(n814), .C(n794), .Z(n812) );
  AO7SVTX6 U482 ( .A(n823), .B(n826), .C(n825), .Z(n816) );
  AO6SVTX6 U483 ( .A(n909), .B(n213), .C(n783), .Z(n826) );
  F_ND2SVTX1 U484 ( .A(n820), .B(n819), .Z(n821) );
  B_ND2SVTX2 U485 ( .A(n829), .B(n828), .Z(n830) );
  B_ND2SVTX2 U486 ( .A(n815), .B(n814), .Z(n817) );
  IVSVTX2 U487 ( .A(n829), .Z(n751) );
  B_ND2SVTX2 U488 ( .A(n782), .B(n781), .Z(n908) );
  IVSVTX2 U489 ( .A(n836), .Z(n747) );
  B_ND2SVTX2 U490 ( .A(n796), .B(n795), .Z(n811) );
  FAS1SVTX2 U491 ( .A(n777), .B(n776), .CI(n775), .CO(n782), .Z(n773) );
  FA1SVTX1 U492 ( .A(n788), .B(n787), .CI(n786), .CO(n793), .Z(n784) );
  B_ND2SVTX2 U493 ( .A(n746), .B(n745), .Z(n834) );
  FA1SVTX4 U494 ( .A(n754), .B(n753), .CI(n752), .CO(n774), .Z(n749) );
  F_ND2ASVTX2 U495 ( .A(n731), .B(n730), .Z(n753) );
  F_ND2SVTX1 U496 ( .A(n760), .B(n211), .Z(n730) );
  AO6SVTX4 U497 ( .A(n849), .B(n847), .C(n554), .Z(n555) );
  AO17SVTX4 U498 ( .A(n682), .B(n681), .C(n685), .D(n680), .Z(n683) );
  B_ND2SVTX1 U499 ( .A(n585), .B(n586), .Z(n565) );
  AO6SVTX4 U500 ( .A(n853), .B(n855), .C(n549), .Z(n842) );
  B_ND2SVTX1 U501 ( .A(n864), .B(n863), .Z(n866) );
  AO6SVTX2 U502 ( .A(n867), .B(n872), .C(n524), .Z(n525) );
  B_ND2SVTX1 U503 ( .A(n677), .B(n584), .Z(n588) );
  B_ND2SVTX1 U504 ( .A(n739), .B(n763), .Z(n740) );
  B_ND2SVTX2 U505 ( .A(n679), .B(n733), .Z(n681) );
  B_ND2SVTX1 U506 ( .A(n848), .B(n847), .Z(n852) );
  B_ND2SVTX1 U507 ( .A(n854), .B(n853), .Z(n857) );
  CTIVSVTX2 U508 ( .A(n868), .Z(n524) );
  B_ND2SVTX1 U509 ( .A(n868), .B(n867), .Z(n874) );
  B_ND2SVTX2 U510 ( .A(n858), .B(n853), .Z(n841) );
  B_ND2SVTX1 U511 ( .A(n567), .B(n566), .Z(n569) );
  CTIVSVTX2 U512 ( .A(n848), .Z(n554) );
  IVSVTX2 U513 ( .A(n567), .Z(n562) );
  B_ND2SVTX2 U514 ( .A(n880), .B(n867), .Z(n526) );
  OR2SVTX2 U515 ( .A(n703), .B(n701), .Z(n761) );
  B_ND2SVTX2 U516 ( .A(n564), .B(n563), .Z(n864) );
  B_ND2SVTX2 U517 ( .A(n523), .B(n522), .Z(n868) );
  B_ND2SVTX2 U518 ( .A(n703), .B(n701), .Z(n762) );
  B_ND2SVTX2 U519 ( .A(n737), .B(n735), .Z(n682) );
  B_ND2SVTX2 U520 ( .A(n561), .B(n560), .Z(n567) );
  B_ND2SVTX1 U521 ( .A(n715), .B(n714), .Z(n723) );
  B_ND2SVTX2 U522 ( .A(n583), .B(n582), .Z(n677) );
  B_ND2SVTX2 U523 ( .A(n551), .B(n550), .Z(n839) );
  B_ND2SVTX2 U524 ( .A(n553), .B(n552), .Z(n848) );
  B_ND2SVTX2 U525 ( .A(n728), .B(n727), .Z(n680) );
  OR2SVTX4 U526 ( .A(n553), .B(n552), .Z(n847) );
  B_ND2SVTX2 U527 ( .A(n548), .B(n547), .Z(n854) );
  B_ND2SVTX2 U528 ( .A(n722), .B(n720), .Z(n739) );
  B_ND2SVTX2 U529 ( .A(n559), .B(n440), .Z(n585) );
  AO7SVTX2 U530 ( .A(n481), .B(n480), .C(n479), .Z(n485) );
  IVSVTX2 U531 ( .A(n881), .Z(n872) );
  B_ND2SVTX1 U532 ( .A(n876), .B(n875), .Z(n879) );
  B_ND2SVTX2 U533 ( .A(n521), .B(n520), .Z(n881) );
  B_ND2SVTX1 U534 ( .A(n905), .B(n904), .Z(n906) );
  B_ND2SVTX1 U535 ( .A(n885), .B(n884), .Z(n887) );
  B_ND2SVTX2 U536 ( .A(n875), .B(n884), .Z(n871) );
  B_ND2SVTX1 U537 ( .A(n900), .B(n899), .Z(n902) );
  EOSVTX2 U538 ( .A(n728), .B(n437), .Z(n581) );
  B_ND2SVTX1 U539 ( .A(n894), .B(n893), .Z(n897) );
  B_ND2SVTX2 U540 ( .A(n517), .B(n516), .Z(n876) );
  B_ND2SVTX2 U541 ( .A(n888), .B(n589), .Z(n513) );
  B_ND2SVTX2 U542 ( .A(n499), .B(n498), .Z(n900) );
  B_ND2SVTX2 U543 ( .A(n488), .B(n487), .Z(n905) );
  B_ND2SVTX2 U544 ( .A(n501), .B(n500), .Z(n894) );
  B_ND2SVTX2 U545 ( .A(n470), .B(n469), .Z(n471) );
  B_ND2SVTX2 U546 ( .A(n508), .B(n507), .Z(n889) );
  B_ND2SVTX2 U547 ( .A(n510), .B(n509), .Z(n590) );
  B_ND2SVTX2 U548 ( .A(n515), .B(n514), .Z(n885) );
  B_ND2SVTX2 U549 ( .A(n450), .B(n435), .Z(n436) );
  ND2SVTX2 U550 ( .A(n403), .B(n402), .Z(n404) );
  IVSVTX4 U551 ( .A(n758), .Z(n445) );
  F_AN2SVTX2 U552 ( .A(n648), .B(n744), .Z(n731) );
  B_ND2SVTX2 U553 ( .A(n620), .B(n619), .Z(n667) );
  IVSVTX2 U554 ( .A(n564), .Z(n529) );
  B_ND2SVTX2 U555 ( .A(n418), .B(n532), .Z(n434) );
  IVSVTX2 U556 ( .A(n553), .Z(n532) );
  AO3SVTX2 U557 ( .A(n641), .B(n633), .C(n632), .D(n631), .Z(n715) );
  B_ND2SVTX2 U558 ( .A(n460), .B(n390), .Z(n455) );
  B_ND2SVTX2 U559 ( .A(n354), .B(n353), .Z(n355) );
  AO7SVTX2 U560 ( .A(O[28]), .B(n597), .C(n289), .Z(n317) );
  NR2SVTX2 U561 ( .A(n623), .B(n633), .Z(n319) );
  AO2SVTX1 U562 ( .A(n636), .B(n422), .C(n630), .D(n413), .Z(n273) );
  B_ND2SVTX1 U563 ( .A(n636), .B(n629), .Z(n613) );
  AO2SVTX1 U564 ( .A(n629), .B(n571), .C(n570), .D(n606), .Z(n574) );
  B_ND2SVTX1 U565 ( .A(n630), .B(n629), .Z(n631) );
  AO4SVTX2 U566 ( .A(n373), .B(n352), .C(n351), .D(n350), .Z(n478) );
  B_ND2SVTX1 U567 ( .A(n637), .B(n636), .Z(n638) );
  CTIVSVTX2 U568 ( .A(n499), .Z(n212) );
  B_ND2SVTX1 U569 ( .A(n606), .B(n630), .Z(n604) );
  IVSVTX2 U570 ( .A(n633), .Z(n636) );
  IVSVTX2 U571 ( .A(n409), .Z(n420) );
  B_ND2SVTX1 U572 ( .A(n637), .B(n630), .Z(n576) );
  IVSVTX2 U573 ( .A(n572), .Z(n351) );
  B_ND2SVTX2 U574 ( .A(O[28]), .B(n274), .Z(n400) );
  B_ND2SVTX2 U575 ( .A(N[0]), .B(O[27]), .Z(n352) );
  NR3SVTX2 U576 ( .A(N[2]), .B(n347), .C(n252), .Z(n230) );
  B_ND2SVTX2 U577 ( .A(n227), .B(n303), .Z(n228) );
  NR4SVTX4 U578 ( .A(N[24]), .B(N[27]), .C(N[26]), .D(N[25]), .Z(n217) );
  NR4SVTX4 U579 ( .A(N[23]), .B(N[21]), .C(N[22]), .D(N[20]), .Z(n246) );
  AO39SVTX2 U580 ( .A(n626), .B(n578), .C(n624), .D(n641), .E(n622), .F(n625), 
        .Z(n333) );
  AO11NSVTX2 U581 ( .A(n488), .B(n719), .C(n717), .D(n212), .E(n672), .F(n463), 
        .Z(n477) );
  EOSVTX8 U582 ( .A(n618), .B(n696), .Z(n729) );
  AO11NSVTX4 U583 ( .A(n722), .B(n689), .C(n445), .D(n686), .E(n672), .F(n674), 
        .Z(n727) );
  EOSVTX4 U584 ( .A(n917), .B(n916), .Z(O[26]) );
  F_IVSVTX0H U585 ( .A(n391), .Z(n393) );
  ND3ABSVTX4 U586 ( .A(n676), .B(n678), .C(n675), .Z(n732) );
  F_ND2SVTX0H U587 ( .A(n645), .B(n669), .Z(n437) );
  AO6SVTX4 U588 ( .A(n528), .B(n869), .C(n527), .Z(n840) );
  NR2SVTX2 U589 ( .A(n551), .B(n550), .Z(n837) );
  AO39SVTX1 U590 ( .A(n626), .B(n623), .C(n624), .D(n621), .E(n622), .F(n602), 
        .Z(n612) );
  AO11NSVTX1 U591 ( .A(n672), .B(n504), .C(n689), .D(n515), .E(n505), .F(n717), 
        .Z(n507) );
  IVSVTX0H U592 ( .A(n840), .Z(n860) );
  AO7SVTX6 U593 ( .A(n840), .B(n556), .C(n555), .Z(n568) );
  NR2SVTX2 U594 ( .A(n583), .B(n582), .Z(n678) );
  AO7SVTX2 U595 ( .A(n744), .B(n771), .C(n743), .Z(n836) );
  IVSVTX0H U596 ( .A(n913), .Z(n699) );
  B_ND2SVTX0H U597 ( .A(N[23]), .B(n572), .Z(n573) );
  IVSVTX2 U598 ( .A(n450), .Z(n537) );
  AO2SVTX1 U599 ( .A(n570), .B(n413), .C(n326), .D(n412), .Z(n328) );
  F_ND2SVTX0H U600 ( .A(n764), .B(n763), .Z(n768) );
  AO7SVTX4 U601 ( .A(n695), .B(n767), .C(n694), .Z(n711) );
  AO2SVTX1 U602 ( .A(N[6]), .B(n306), .C(n363), .D(N[22]), .Z(n307) );
  IVSVTX6 U603 ( .A(n248), .Z(n359) );
  AO2SVTX1 U604 ( .A(n253), .B(n225), .C(N[13]), .D(n315), .Z(n226) );
  EOSVTX0H U605 ( .A(n907), .B(n906), .Z(O[0]) );
  EOSVTX0H U606 ( .A(n902), .B(n901), .Z(O[1]) );
  ENSVTX0H U607 ( .A(n897), .B(n896), .Z(O[2]) );
  ENSVTX0H U608 ( .A(n891), .B(n890), .Z(O[3]) );
  EOSVTX0H U609 ( .A(n594), .B(n593), .Z(O[4]) );
  EOSVTX0H U610 ( .A(n887), .B(n886), .Z(O[5]) );
  ENSVTX0H U611 ( .A(n879), .B(n878), .Z(O[6]) );
  ENSVTX0H U612 ( .A(n883), .B(n882), .Z(O[7]) );
  ENSVTX0H U613 ( .A(n861), .B(n860), .Z(O[9]) );
  EOSVTX0H U614 ( .A(n857), .B(n856), .Z(O[10]) );
  AO6SVTX1 U615 ( .A(n860), .B(n858), .C(n855), .Z(n856) );
  EOSVTX0H U616 ( .A(n846), .B(n845), .Z(O[11]) );
  EOSVTX0H U617 ( .A(n852), .B(n851), .Z(O[12]) );
  EOSVTX0H U618 ( .A(n866), .B(n865), .Z(O[14]) );
  EOSVTX0H U619 ( .A(n588), .B(n587), .Z(O[16]) );
  AO6CSVTX1 U620 ( .A(n675), .B(n586), .C(n585), .Z(n587) );
  ENSVTX0H U621 ( .A(n836), .B(n835), .Z(O[17]) );
  EOSVTX0H U622 ( .A(n914), .B(n913), .Z(n917) );
  IVSVTX0H U623 ( .A(n463), .Z(n488) );
  OR2SVTX2 U624 ( .A(n782), .B(n781), .Z(n213) );
  FA1SVTX1 U625 ( .A(n802), .B(n801), .CI(1'b0), .CO(n803), .Z(n795) );
  IVSVTX4 U626 ( .A(n264), .Z(n325) );
  IVSVTX6 U627 ( .A(n325), .Z(n363) );
  IVSVTX2 U628 ( .A(n263), .Z(n281) );
  IVSVTX2 U629 ( .A(n344), .Z(n373) );
  OR2SVTX2 U630 ( .A(n700), .B(n699), .Z(n214) );
  NR2SVTX2 U631 ( .A(N[28]), .B(N[31]), .Z(n216) );
  NR2SVTX2 U632 ( .A(N[30]), .B(N[29]), .Z(n215) );
  ND2SVTX4 U633 ( .A(n216), .B(n215), .Z(n248) );
  IVSVTX0H U634 ( .A(N[26]), .Z(n220) );
  IVSVTX0H U635 ( .A(N[29]), .Z(n218) );
  AO8SVTX1 U636 ( .A(N[25]), .B(n220), .C(n359), .D(n219), .Z(n221) );
  IVSVTX2 U637 ( .A(N[18]), .Z(n303) );
  NR2ASVTX6 U638 ( .A(n246), .B(n260), .Z(n231) );
  NR3ABSVTX2 U639 ( .A(N[17]), .B(n303), .C(n251), .Z(n240) );
  NR4SVTX2 U640 ( .A(N[4]), .B(N[5]), .C(N[6]), .D(N[7]), .Z(n242) );
  NR2SVTX2 U641 ( .A(N[11]), .B(N[9]), .Z(n224) );
  NR2SVTX2 U642 ( .A(N[8]), .B(N[10]), .Z(n223) );
  IVSVTX2 U643 ( .A(N[15]), .Z(n267) );
  NR2SVTX2 U644 ( .A(N[13]), .B(N[12]), .Z(n222) );
  ND3SVTX4 U645 ( .A(n267), .B(n315), .C(n222), .Z(n243) );
  NR3ABSVTX2 U646 ( .A(n224), .B(n223), .C(n243), .Z(n245) );
  ND2SVTX4 U647 ( .A(n242), .B(n245), .Z(n252) );
  IVSVTX4 U648 ( .A(n245), .Z(n262) );
  IVSVTX2 U649 ( .A(n243), .Z(n253) );
  NR2SVTX2 U650 ( .A(N[10]), .B(n286), .Z(n225) );
  ND4ABCSVTX8 U651 ( .A(N[17]), .B(N[19]), .C(n228), .D(n231), .Z(O[31]) );
  IVSVTX2 U652 ( .A(O[31]), .Z(n301) );
  AO7SVTX2 U653 ( .A(n230), .B(n229), .C(n301), .Z(n239) );
  NR2ASVTX1 U654 ( .A(N[23]), .B(n260), .Z(n232) );
  IVSVTX0H U655 ( .A(N[7]), .Z(n358) );
  AO6SVTX2 U656 ( .A(n253), .B(N[11]), .C(N[15]), .Z(n233) );
  AO7SVTX4 U657 ( .A(n358), .B(n262), .C(n233), .Z(n235) );
  NR2ASVTX2 U658 ( .A(N[3]), .B(n252), .Z(n234) );
  AO6ABSVTX2 U659 ( .A(n235), .B(n234), .C(O[31]), .Z(n236) );
  ND4ABSVTX8 U660 ( .A(n241), .B(n240), .C(n239), .D(n389), .Z(O[27]) );
  IVSVTX0H U661 ( .A(n242), .Z(n244) );
  NR2SVTX2 U662 ( .A(n246), .B(n260), .Z(n247) );
  AO3CDSVTX4 U663 ( .A(O[31]), .B(n249), .C(n248), .D(n247), .Z(O[29]) );
  IVSVTX4 U664 ( .A(O[29]), .Z(n366) );
  AO6SVTX1 U665 ( .A(n359), .B(N[26]), .C(N[30]), .Z(n250) );
  NR2ASVTX2 U666 ( .A(N[18]), .B(n251), .Z(n258) );
  IVSVTX0H U667 ( .A(n252), .Z(n256) );
  AO6SVTX1 U668 ( .A(n253), .B(N[10]), .C(N[14]), .Z(n254) );
  AO7SVTX1 U669 ( .A(n360), .B(n262), .C(n254), .Z(n255) );
  AO17SVTX2 U670 ( .A(n256), .B(N[2]), .C(n255), .D(n301), .Z(n257) );
  ND4ABSVTX8 U671 ( .A(n259), .B(n258), .C(n257), .D(n389), .Z(O[28]) );
  AN2SVTX4 U672 ( .A(O[27]), .B(n326), .Z(n630) );
  IVSVTX2 U673 ( .A(n260), .Z(n261) );
  ND2SVTX4 U674 ( .A(O[31]), .B(n263), .Z(n343) );
  IVSVTX4 U675 ( .A(n343), .Z(n384) );
  NR2ASVTX2 U676 ( .A(O[31]), .B(n263), .Z(n264) );
  AO2SVTX2 U677 ( .A(n384), .B(N[13]), .C(n363), .D(N[5]), .Z(n410) );
  AO2SVTX2 U678 ( .A(n384), .B(N[12]), .C(n363), .D(N[4]), .Z(n406) );
  AO4SVTX1 U679 ( .A(n640), .B(n410), .C(n406), .D(n633), .Z(n270) );
  IVSVTX4 U680 ( .A(n281), .Z(O[30]) );
  F_ND2ASVTX2 U681 ( .A(O[31]), .B(O[30]), .Z(n312) );
  IVSVTX4 U682 ( .A(n312), .Z(n305) );
  AO11SVTX4 U683 ( .A(N[18]), .B(n384), .C(n363), .D(N[10]), .E(n305), .F(N[2]), .Z(n641) );
  AO4SVTX1 U684 ( .A(n325), .B(n360), .C(n343), .D(n315), .Z(n422) );
  AO11SVTX4 U685 ( .A(n384), .B(N[16]), .C(n363), .D(N[8]), .E(n305), .F(N[0]), 
        .Z(n578) );
  IVSVTX2 U686 ( .A(n578), .Z(n265) );
  AO11SVTX2 U687 ( .A(n266), .B(n421), .C(n422), .D(n571), .E(n265), .F(n570), 
        .Z(n323) );
  AO11NSVTX2 U688 ( .A(N[3]), .B(n305), .C(N[19]), .D(n384), .E(n363), .F(
        N[11]), .Z(n629) );
  AO4SVTX1 U689 ( .A(n325), .B(n358), .C(n267), .D(n343), .Z(n413) );
  IVSVTX0H U690 ( .A(N[17]), .Z(n268) );
  AO39SVTX2 U691 ( .A(n268), .B(n343), .C(n347), .D(n312), .E(n325), .F(n286), 
        .Z(n637) );
  AO11SVTX2 U692 ( .A(n629), .B(n421), .C(n413), .D(n571), .E(n637), .F(n570), 
        .Z(n332) );
  F_MUX21NSVTX0H U693 ( .A(n323), .B(n332), .S(O[27]), .Z(n269) );
  OR2SVTX2 U694 ( .A(n270), .B(n269), .Z(n559) );
  AO11SVTX2 U695 ( .A(n384), .B(N[20]), .C(n363), .D(N[12]), .E(n305), .F(N[4]), .Z(n625) );
  IVSVTX0H U696 ( .A(N[13]), .Z(n284) );
  AO39SVTX2 U697 ( .A(n271), .B(n343), .C(n365), .D(n312), .E(n284), .F(n325), 
        .Z(n606) );
  AO11NSVTX4 U698 ( .A(n637), .B(n571), .C(n629), .D(n570), .E(n606), .F(n421), 
        .Z(n320) );
  ND2SVTX2 U699 ( .A(n273), .B(n272), .Z(n737) );
  NR2SVTX2 U700 ( .A(O[29]), .B(n343), .Z(n387) );
  IVSVTX0H U701 ( .A(N[19]), .Z(n276) );
  AO6SVTX1 U702 ( .A(n301), .B(N[11]), .C(N[27]), .Z(n275) );
  AO7SVTX1 U703 ( .A(n276), .B(O[30]), .C(n275), .Z(n277) );
  AO6SVTX1 U704 ( .A(N[3]), .B(n306), .C(n277), .Z(n278) );
  AO2SVTX4 U705 ( .A(n305), .B(N[7]), .C(n363), .D(N[15]), .Z(n607) );
  F_MUX21NSVTX1 U706 ( .A(n278), .B(n607), .S(n366), .Z(n279) );
  NR2ASVTX1 U707 ( .A(n280), .B(n279), .Z(n597) );
  AO6SVTX1 U708 ( .A(n281), .B(N[21]), .C(N[29]), .Z(n282) );
  AO3SVTX1 U709 ( .A(n312), .B(n284), .C(n283), .D(n282), .Z(n288) );
  NR2ASVTX1 U710 ( .A(N[17]), .B(n263), .Z(n285) );
  AO1ABSVTX1 U711 ( .A(O[31]), .B(n286), .C(N[25]), .D(n285), .Z(n287) );
  AO7SVTX2 U712 ( .A(n298), .B(n347), .C(n287), .Z(n595) );
  IVSVTX0H U713 ( .A(N[8]), .Z(n291) );
  IVSVTX0H U714 ( .A(N[24]), .Z(n290) );
  AO7SVTX1 U715 ( .A(n291), .B(O[31]), .C(n290), .Z(n294) );
  NR2ASVTX1 U716 ( .A(N[16]), .B(n263), .Z(n293) );
  ND3ABSVTX2 U717 ( .A(n294), .B(n293), .C(n292), .Z(n601) );
  IVSVTX0H U718 ( .A(N[20]), .Z(n296) );
  IVSVTX0H U719 ( .A(N[28]), .Z(n295) );
  AO7SVTX1 U720 ( .A(n296), .B(n325), .C(n295), .Z(n300) );
  IVSVTX0H U721 ( .A(N[4]), .Z(n357) );
  IVSVTX0H U722 ( .A(N[12]), .Z(n297) );
  AO4SVTX1 U723 ( .A(n298), .B(n357), .C(n312), .D(n297), .Z(n299) );
  NR2SVTX2 U724 ( .A(O[28]), .B(n316), .Z(n310) );
  IVSVTX0H U725 ( .A(N[2]), .Z(n361) );
  AO6SVTX1 U726 ( .A(n301), .B(N[10]), .C(N[26]), .Z(n302) );
  AO7SVTX1 U727 ( .A(n303), .B(n263), .C(n302), .Z(n304) );
  AO6SVTX1 U728 ( .A(n305), .B(N[14]), .C(N[30]), .Z(n308) );
  AO3SVTX1 U729 ( .A(n602), .B(n626), .C(n308), .D(n307), .Z(n309) );
  AO2ABSVTX4 U730 ( .C(n274), .D(n311), .A(n310), .B(n309), .Z(n760) );
  AO4SVTX1 U731 ( .A(n343), .B(n313), .C(n360), .D(n312), .Z(n314) );
  AO6ABSVTX2 U732 ( .A(n315), .B(n325), .C(n314), .Z(n623) );
  AO4SVTX1 U733 ( .A(n316), .B(n596), .C(n602), .D(n624), .Z(n598) );
  OR2SVTX2 U734 ( .A(n760), .B(n648), .Z(n911) );
  IVSVTX2 U735 ( .A(n648), .Z(n698) );
  ND2SVTX4 U736 ( .A(n760), .B(n698), .Z(n758) );
  AO39SVTX1 U737 ( .A(n626), .B(n641), .C(n624), .D(n625), .E(n622), .F(n623), 
        .Z(n575) );
  AO3SVTX4 U738 ( .A(n578), .B(n640), .C(n322), .D(n321), .Z(n728) );
  IVSVTX0H U739 ( .A(n323), .Z(n329) );
  IVSVTX0H U740 ( .A(N[3]), .Z(n374) );
  IVSVTX0H U741 ( .A(N[11]), .Z(n324) );
  AO4SVTX1 U742 ( .A(n325), .B(n374), .C(n324), .D(n343), .Z(n412) );
  AO3SVTX2 U743 ( .A(n410), .B(n626), .C(n328), .D(n327), .Z(n407) );
  F_MUX21NSVTX1 U744 ( .A(n329), .B(n407), .S(n274), .Z(n330) );
  AO7SVTX2 U745 ( .A(n406), .B(n640), .C(n330), .Z(n564) );
  IVSVTX0H U746 ( .A(n737), .Z(n338) );
  F_IVSVTX0H U747 ( .A(n332), .Z(n334) );
  AO3SVTX2 U748 ( .A(n410), .B(n633), .C(n336), .D(n335), .Z(n583) );
  IVSVTX0H U749 ( .A(n583), .Z(n337) );
  ND2SVTX2 U750 ( .A(n338), .B(n337), .Z(n339) );
  NR2SVTX2 U751 ( .A(n441), .B(n339), .Z(n645) );
  IVSVTX4 U752 ( .A(n387), .Z(n364) );
  IVSVTX0H U753 ( .A(N[0]), .Z(n340) );
  IVSVTX0H U754 ( .A(n375), .Z(n342) );
  NR2ASVTX2 U755 ( .A(n384), .B(n622), .Z(n572) );
  AO7SVTX1 U756 ( .A(n389), .B(n342), .C(n341), .Z(n346) );
  NR2SVTX2 U757 ( .A(n624), .B(n343), .Z(n344) );
  NR2SVTX0H U758 ( .A(n350), .B(n373), .Z(n345) );
  NR2SVTX2 U759 ( .A(n346), .B(n345), .Z(n463) );
  AO4SVTX1 U760 ( .A(n364), .B(n347), .C(n365), .D(n359), .Z(n362) );
  MUX21NSVTX2 U761 ( .A(n375), .B(n362), .S(O[27]), .Z(n372) );
  F_MUX21NSVTX1 U762 ( .A(N[2]), .B(N[3]), .S(O[27]), .Z(n348) );
  AO4SVTX2 U763 ( .A(n372), .B(n596), .C(n348), .D(n373), .Z(n499) );
  NR2SVTX2 U764 ( .A(n352), .B(n351), .Z(n470) );
  NR2SVTX2 U765 ( .A(n473), .B(n470), .Z(n354) );
  AO4SVTX2 U766 ( .A(n373), .B(n349), .C(n351), .D(n348), .Z(n483) );
  NR2SVTX2 U767 ( .A(n483), .B(n478), .Z(n353) );
  NR2SVTX2 U768 ( .A(n356), .B(n355), .Z(n464) );
  AO2SVTX2 U769 ( .A(n384), .B(N[8]), .C(n363), .D(N[0]), .Z(n426) );
  AO4SVTX2 U770 ( .A(n426), .B(n366), .C(n357), .D(n364), .Z(n367) );
  AO4SVTX1 U771 ( .A(n364), .B(n374), .C(n358), .D(n359), .Z(n369) );
  MUX21NSVTX2 U772 ( .A(n367), .B(n369), .S(n274), .Z(n385) );
  AO4SVTX1 U773 ( .A(n364), .B(n361), .C(n360), .D(n359), .Z(n368) );
  AO2SVTX2 U774 ( .A(n384), .B(N[9]), .C(n363), .D(N[1]), .Z(n427) );
  AO4SVTX1 U775 ( .A(n427), .B(n366), .C(n365), .D(n364), .Z(n396) );
  MUX21NSVTX2 U776 ( .A(n396), .B(n367), .S(n274), .Z(n388) );
  F_MUX21NSVTX1 U777 ( .A(n369), .B(n368), .S(n274), .Z(n371) );
  MUX21NSVTX2 U778 ( .A(n388), .B(n371), .S(n596), .Z(n515) );
  IVSVTX0H U779 ( .A(n515), .Z(n370) );
  ND2SVTX2 U780 ( .A(n493), .B(n370), .Z(n382) );
  MUX21NSVTX2 U781 ( .A(n372), .B(n371), .S(O[28]), .Z(n508) );
  IVSVTX0H U782 ( .A(n508), .Z(n381) );
  NR2ASVTX1 U783 ( .A(n375), .B(O[28]), .Z(n376) );
  IVSVTX2 U784 ( .A(n501), .Z(n380) );
  ND2SVTX2 U785 ( .A(n381), .B(n380), .Z(n491) );
  NR2SVTX2 U786 ( .A(n382), .B(n491), .Z(n383) );
  ND2SVTX4 U787 ( .A(n464), .B(n383), .Z(n447) );
  IVSVTX0H U788 ( .A(n396), .Z(n386) );
  AO2SVTX2 U789 ( .A(n420), .B(O[29]), .C(N[6]), .D(n387), .Z(n391) );
  AO39SVTX2 U790 ( .A(n400), .B(n386), .C(n389), .D(n391), .E(O[28]), .F(n385), 
        .Z(n517) );
  IVSVTX2 U791 ( .A(n517), .Z(n460) );
  AO2SVTX2 U792 ( .A(n412), .B(O[29]), .C(N[7]), .D(n387), .Z(n401) );
  AO39SVTX2 U793 ( .A(n389), .B(n401), .C(n400), .D(n391), .E(O[28]), .F(n388), 
        .Z(n521) );
  IVSVTX2 U794 ( .A(n406), .Z(n419) );
  IVSVTX0H U795 ( .A(n426), .Z(n392) );
  AO11SVTX2 U796 ( .A(n393), .B(n596), .C(n419), .D(n421), .E(n392), .F(n571), 
        .Z(n395) );
  AO39SVTX1 U797 ( .A(n622), .B(n410), .C(n626), .D(n427), .E(O[28]), .F(n401), 
        .Z(n423) );
  MUX21NSVTX2 U798 ( .A(n395), .B(n394), .S(O[27]), .Z(n546) );
  IVSVTX2 U799 ( .A(n546), .Z(n403) );
  IVSVTX2 U800 ( .A(n395), .Z(n398) );
  NR2ASVTX1 U801 ( .A(n396), .B(O[28]), .Z(n397) );
  IVSVTX2 U802 ( .A(n523), .Z(n402) );
  NR2SVTX2 U803 ( .A(n455), .B(n404), .Z(n450) );
  IVSVTX0H U804 ( .A(n422), .Z(n405) );
  AO39SVTX2 U805 ( .A(n626), .B(n406), .C(n624), .D(n405), .E(n622), .F(n578), 
        .Z(n414) );
  MUX21NSVTX2 U806 ( .A(n407), .B(n414), .S(n274), .Z(n408) );
  AO7SVTX2 U807 ( .A(n409), .B(n633), .C(n408), .Z(n561) );
  IVSVTX0H U808 ( .A(n410), .Z(n411) );
  AO11SVTX2 U809 ( .A(n413), .B(n421), .C(n412), .D(n571), .E(n411), .F(n570), 
        .Z(n429) );
  MUX21NSVTX2 U810 ( .A(n415), .B(n414), .S(O[27]), .Z(n417) );
  AO3SVTX4 U811 ( .A(n427), .B(n633), .C(n417), .D(n416), .Z(n553) );
  AO11SVTX2 U812 ( .A(n422), .B(n421), .C(n420), .D(n571), .E(n419), .F(n570), 
        .Z(n428) );
  IVSVTX0H U813 ( .A(n428), .Z(n424) );
  MUX21NSVTX2 U814 ( .A(n424), .B(n423), .S(n274), .Z(n425) );
  AO7SVTX4 U815 ( .A(n426), .B(n640), .C(n425), .Z(n548) );
  IVSVTX2 U816 ( .A(n548), .Z(n433) );
  AO4SVTX1 U817 ( .A(n640), .B(n427), .C(n426), .D(n633), .Z(n431) );
  F_MUX21NSVTX1 U818 ( .A(n429), .B(n428), .S(n274), .Z(n430) );
  NR2SVTX2 U819 ( .A(n434), .B(n538), .Z(n435) );
  AN2ABSVTX8 U820 ( .A(n447), .B(n436), .Z(n669) );
  NR2SVTX0H U821 ( .A(n583), .B(n441), .Z(n438) );
  ND2SVTX2 U822 ( .A(n438), .B(n669), .Z(n439) );
  AO11NSVTX2 U823 ( .A(n737), .B(n689), .C(n445), .D(n581), .E(n687), .F(n444), 
        .Z(n440) );
  NR2SVTX2 U824 ( .A(n559), .B(n440), .Z(n676) );
  IVSVTX0H U825 ( .A(n676), .Z(n586) );
  IVSVTX0H U826 ( .A(n441), .Z(n442) );
  EOSVTX0H U827 ( .A(n583), .B(n443), .Z(n558) );
  AO11NSVTX1 U828 ( .A(n583), .B(n689), .C(n445), .D(n444), .E(n687), .F(n558), 
        .Z(n563) );
  NR2SVTX2 U829 ( .A(n564), .B(n563), .Z(n862) );
  EOSVTX2 U830 ( .A(n548), .B(n446), .Z(n453) );
  OR2SVTX2 U831 ( .A(n523), .B(n455), .Z(n448) );
  NR2SVTX2 U832 ( .A(n448), .B(n447), .Z(n449) );
  ENSVTX0H U833 ( .A(n546), .B(n449), .Z(n454) );
  AO11NSVTX2 U834 ( .A(n546), .B(n719), .C(n717), .D(n453), .E(n672), .F(n454), 
        .Z(n520) );
  OR2SVTX2 U835 ( .A(n521), .B(n520), .Z(n880) );
  NR2SVTX2 U836 ( .A(n548), .B(n537), .Z(n451) );
  AO11NSVTX4 U837 ( .A(n548), .B(n719), .C(n717), .D(n542), .E(n672), .F(n453), 
        .Z(n522) );
  OR2SVTX4 U838 ( .A(n523), .B(n522), .Z(n867) );
  F_AO2SVTX1 U839 ( .A(n454), .B(n717), .C(n719), .D(n523), .Z(n459) );
  IVSVTX0H U840 ( .A(n455), .Z(n456) );
  F_EOSVTX2 U841 ( .A(n523), .B(n457), .Z(n462) );
  ND2SVTX2 U842 ( .A(n459), .B(n458), .Z(n516) );
  OR2SVTX2 U843 ( .A(n517), .B(n516), .Z(n875) );
  ND2SVTX2 U844 ( .A(n460), .B(n540), .Z(n461) );
  AO11NSVTX2 U845 ( .A(n521), .B(n719), .C(n717), .D(n462), .E(n672), .F(n506), 
        .Z(n514) );
  NR2SVTX2 U846 ( .A(n515), .B(n514), .Z(n877) );
  NR2SVTX2 U847 ( .A(n526), .B(n871), .Z(n528) );
  NR2SVTX2 U848 ( .A(n501), .B(n495), .Z(n465) );
  ENSVTX0H U849 ( .A(n508), .B(n465), .Z(n490) );
  F_EOSVTX2 U850 ( .A(n501), .B(n495), .Z(n466) );
  NR2SVTX2 U851 ( .A(n488), .B(n487), .Z(n903) );
  AO11NSVTX1 U852 ( .A(n499), .B(n719), .C(n717), .D(n466), .E(n672), .F(n212), 
        .Z(n482) );
  OR2SVTX2 U853 ( .A(n483), .B(n482), .Z(n486) );
  NR2SVTX2 U854 ( .A(n478), .B(n477), .Z(n481) );
  IVSVTX0H U855 ( .A(n483), .Z(n468) );
  AO11NSVTX4 U856 ( .A(n483), .B(n719), .C(n717), .D(n463), .E(n672), .F(n468), 
        .Z(n472) );
  OR2SVTX2 U857 ( .A(n473), .B(n472), .Z(n476) );
  IVSVTX0H U858 ( .A(n478), .Z(n467) );
  AO11NSVTX2 U859 ( .A(n478), .B(n719), .C(n717), .D(n468), .E(n672), .F(n467), 
        .Z(n469) );
  F_IVSVTX0H U860 ( .A(n471), .Z(n475) );
  F_AN2SVTX2 U861 ( .A(n473), .B(n472), .Z(n474) );
  AO6SVTX2 U862 ( .A(n476), .B(n475), .C(n474), .Z(n480) );
  F_AN2SVTX2 U863 ( .A(n483), .B(n482), .Z(n484) );
  NR2SVTX2 U864 ( .A(n491), .B(n495), .Z(n489) );
  ENSVTX0H U865 ( .A(n510), .B(n489), .Z(n497) );
  NR2SVTX2 U866 ( .A(n499), .B(n498), .Z(n898) );
  IVSVTX0H U867 ( .A(n491), .Z(n492) );
  NR2SVTX2 U868 ( .A(n495), .B(n494), .Z(n496) );
  ENSVTX0H U869 ( .A(n515), .B(n496), .Z(n504) );
  AO11NSVTX4 U870 ( .A(n672), .B(n497), .C(n689), .D(n510), .E(n717), .F(n504), 
        .Z(n500) );
  NR2SVTX2 U871 ( .A(n501), .B(n500), .Z(n892) );
  NR2SVTX2 U872 ( .A(n898), .B(n892), .Z(n503) );
  AO7SVTX2 U873 ( .A(n900), .B(n892), .C(n894), .Z(n502) );
  ENSVTX0H U874 ( .A(n517), .B(n540), .Z(n505) );
  OR2SVTX2 U875 ( .A(n508), .B(n507), .Z(n888) );
  AO11NSVTX2 U876 ( .A(n517), .B(n719), .C(n717), .D(n506), .E(n672), .F(n505), 
        .Z(n509) );
  OR2SVTX2 U877 ( .A(n510), .B(n509), .Z(n589) );
  IVSVTX2 U878 ( .A(n889), .Z(n592) );
  IVSVTX0H U879 ( .A(n590), .Z(n511) );
  AO6SVTX2 U880 ( .A(n589), .B(n592), .C(n511), .Z(n512) );
  AO7SVTX4 U881 ( .A(n591), .B(n513), .C(n512), .Z(n869) );
  F_IVSVTX0H U882 ( .A(n885), .Z(n519) );
  IVSVTX0H U883 ( .A(n876), .Z(n518) );
  AO6SVTX2 U884 ( .A(n875), .B(n519), .C(n518), .Z(n870) );
  AO11NSVTX4 U885 ( .A(n564), .B(n719), .C(n445), .D(n557), .E(n687), .F(n536), 
        .Z(n552) );
  IVSVTX1 U886 ( .A(n538), .Z(n531) );
  ND2SVTX2 U887 ( .A(n532), .B(n531), .Z(n533) );
  NR2SVTX2 U888 ( .A(n537), .B(n533), .Z(n534) );
  ND2SVTX2 U889 ( .A(n540), .B(n534), .Z(n535) );
  EOSVTX2 U890 ( .A(n561), .B(n535), .Z(n544) );
  AO11NSVTX2 U891 ( .A(n561), .B(n719), .C(n445), .D(n536), .E(n672), .F(n544), 
        .Z(n550) );
  NR2SVTX2 U892 ( .A(n538), .B(n537), .Z(n539) );
  ND2SVTX2 U893 ( .A(n540), .B(n539), .Z(n541) );
  F_EOSVTX2 U894 ( .A(n553), .B(n541), .Z(n543) );
  AO11NSVTX2 U895 ( .A(n551), .B(n719), .C(n717), .D(n543), .E(n672), .F(n542), 
        .Z(n545) );
  OR2SVTX2 U896 ( .A(n546), .B(n545), .Z(n858) );
  AO11NSVTX2 U897 ( .A(n553), .B(n719), .C(n717), .D(n544), .E(n672), .F(n543), 
        .Z(n547) );
  OR2SVTX4 U898 ( .A(n548), .B(n547), .Z(n853) );
  NR2SVTX2 U899 ( .A(n837), .B(n841), .Z(n850) );
  IVSVTX2 U900 ( .A(n859), .Z(n855) );
  IVSVTX2 U901 ( .A(n854), .Z(n549) );
  AO7SVTX4 U902 ( .A(n837), .B(n842), .C(n839), .Z(n849) );
  AO11NSVTX2 U903 ( .A(n559), .B(n689), .C(n445), .D(n558), .E(n687), .F(n557), 
        .Z(n560) );
  OR2SVTX2 U904 ( .A(n561), .B(n560), .Z(n566) );
  AO6SVTX8 U905 ( .A(n568), .B(n566), .C(n562), .Z(n865) );
  AO7SVTX8 U906 ( .A(n862), .B(n865), .C(n864), .Z(n675) );
  ENSVTX0H U907 ( .A(n565), .B(n675), .Z(O[15]) );
  ENSVTX0H U908 ( .A(n569), .B(n568), .Z(O[13]) );
  AO3SVTX1 U909 ( .A(n607), .B(n622), .C(n574), .D(n573), .Z(n635) );
  F_MUX21NSVTX0H U910 ( .A(n635), .B(n575), .S(n274), .Z(n577) );
  AO3SVTX2 U911 ( .A(n578), .B(n633), .C(n577), .D(n576), .Z(n757) );
  IVSVTX2 U912 ( .A(n645), .Z(n668) );
  NR2SVTX2 U913 ( .A(n728), .B(n668), .Z(n579) );
  ND2SVTX2 U914 ( .A(n579), .B(n669), .Z(n580) );
  AO11NSVTX2 U915 ( .A(n728), .B(n689), .C(n717), .D(n673), .E(n687), .F(n581), 
        .Z(n582) );
  IVSVTX0H U916 ( .A(n678), .Z(n584) );
  IVSVTX0H U917 ( .A(n591), .Z(n890) );
  AO6SVTX1 U918 ( .A(n890), .B(n888), .C(n592), .Z(n593) );
  IVSVTX0H U919 ( .A(n595), .Z(n608) );
  AO4SVTX1 U920 ( .A(n597), .B(n596), .C(n608), .D(n624), .Z(n603) );
  IVSVTX0H U921 ( .A(n601), .Z(n621) );
  IVSVTX0H U922 ( .A(n706), .Z(n616) );
  IVSVTX0H U923 ( .A(n606), .Z(n611) );
  AO4SVTX1 U924 ( .A(n608), .B(n622), .C(n607), .D(n624), .Z(n609) );
  AO6SVTX1 U925 ( .A(N[23]), .B(n344), .C(n609), .Z(n610) );
  AO7SVTX1 U926 ( .A(n611), .B(n626), .C(n610), .Z(n628) );
  AO3SVTX2 U927 ( .A(n625), .B(n640), .C(n614), .D(n613), .Z(n703) );
  IVSVTX0H U928 ( .A(n703), .Z(n615) );
  ND2SVTX2 U929 ( .A(n616), .B(n615), .Z(n651) );
  IVSVTX0H U930 ( .A(n651), .Z(n617) );
  IVSVTX0H U931 ( .A(n728), .Z(n620) );
  AO39SVTX1 U932 ( .A(n626), .B(n625), .C(n624), .D(n623), .E(n622), .F(n621), 
        .Z(n634) );
  IVSVTX0H U933 ( .A(n715), .Z(n642) );
  F_MUX21NSVTX0H U934 ( .A(n635), .B(n634), .S(O[27]), .Z(n639) );
  AO3SVTX2 U935 ( .A(n641), .B(n640), .C(n639), .D(n638), .Z(n722) );
  NR2SVTX2 U936 ( .A(n667), .B(n643), .Z(n644) );
  NR2SVTX2 U937 ( .A(n646), .B(n656), .Z(n647) );
  NR2SVTX2 U938 ( .A(n651), .B(n656), .Z(n652) );
  NR2SVTX2 U939 ( .A(n703), .B(n656), .Z(n654) );
  AO11NSVTX4 U940 ( .A(n706), .B(n689), .C(n445), .D(n660), .E(n687), .F(n659), 
        .Z(n714) );
  NR2SVTX2 U941 ( .A(n715), .B(n714), .Z(n693) );
  IVSVTX0H U942 ( .A(n656), .Z(n657) );
  ND2SVTX2 U943 ( .A(n669), .B(n657), .Z(n658) );
  EOSVTX1 U944 ( .A(n703), .B(n658), .Z(n688) );
  AO11NSVTX4 U945 ( .A(n703), .B(n689), .C(n445), .D(n659), .E(n687), .F(n688), 
        .Z(n720) );
  NR2SVTX2 U946 ( .A(n722), .B(n720), .Z(n738) );
  IVSVTX2 U947 ( .A(n738), .Z(n763) );
  AO11NSVTX4 U948 ( .A(n799), .B(n719), .C(n717), .D(n661), .E(n672), .F(n660), 
        .Z(n701) );
  ND3SVTX2 U949 ( .A(n764), .B(n763), .C(n761), .Z(n695) );
  IVSVTX0H U950 ( .A(n667), .Z(n662) );
  NR2SVTX2 U951 ( .A(n668), .B(n664), .Z(n665) );
  NR2SVTX2 U952 ( .A(n668), .B(n667), .Z(n670) );
  F_EOSVTX2 U953 ( .A(n722), .B(n671), .Z(n674) );
  NR2SVTX2 U954 ( .A(n728), .B(n727), .Z(n685) );
  AO11NSVTX4 U955 ( .A(n757), .B(n689), .C(n445), .D(n674), .E(n687), .F(n673), 
        .Z(n735) );
  NR2SVTX2 U956 ( .A(n737), .B(n735), .Z(n684) );
  IVSVTX0H U957 ( .A(n684), .Z(n679) );
  AO21DSVTX8 U958 ( .A(n685), .B(n684), .C(n732), .D(n683), .Z(n692) );
  OR2SVTX2 U959 ( .A(n757), .B(n755), .Z(n691) );
  F_AN2SVTX2 U960 ( .A(n757), .B(n755), .Z(n690) );
  AO6SVTX8 U961 ( .A(n692), .B(n691), .C(n690), .Z(n767) );
  AO7SVTX2 U962 ( .A(n739), .B(n693), .C(n723), .Z(n765) );
  AO6CSVTX2 U963 ( .A(n765), .B(n761), .C(n762), .Z(n694) );
  AN2ABSVTX6 U964 ( .A(n729), .B(n697), .Z(n789) );
  NR2SVTX2 U965 ( .A(n912), .B(n729), .Z(n716) );
  F_FA1SVTX1 U966 ( .A(n703), .B(n702), .CI(n701), .CO(n705), .Z(n791) );
  AO7SVTX1 U967 ( .A(n709), .B(n211), .C(n707), .Z(n801) );
  NR2SVTX2 U969 ( .A(n796), .B(n795), .Z(n809) );
  AO3SVTX4 U970 ( .A(n771), .B(n709), .C(n708), .D(n758), .Z(n779) );
  IVSVTX0H U971 ( .A(n710), .Z(n712) );
  ENSVTX0H U972 ( .A(n712), .B(n711), .Z(n713) );
  NR2ASVTX2 U973 ( .A(n713), .B(n771), .Z(n778) );
  HA1SVTX1 U974 ( .A(n715), .B(n714), .CO(n702), .S(n788) );
  AO20SVTX2 U975 ( .A(n731), .B(n717), .C(n729), .D(n716), .Z(n718) );
  F_FA1SVTX1 U976 ( .A(n722), .B(n721), .CI(n720), .CO(n786), .Z(n780) );
  AO7SVTX1 U977 ( .A(n738), .B(n767), .C(n739), .Z(n724) );
  ENSVTX0H U978 ( .A(n725), .B(n724), .Z(n726) );
  NR2ASVTX2 U979 ( .A(n726), .B(n771), .Z(n748) );
  HA1SVTX1 U980 ( .A(n728), .B(n727), .CO(n756), .S(n754) );
  NR2SVTX2 U981 ( .A(n748), .B(n749), .Z(n734) );
  IVSVTX2 U982 ( .A(n734), .Z(n828) );
  F_FA1SVTX1 U983 ( .A(n737), .B(n736), .CI(n735), .CO(n752), .Z(n746) );
  NR2SVTX2 U984 ( .A(n746), .B(n745), .Z(n832) );
  AO7SVTX4 U985 ( .A(n832), .B(n747), .C(n834), .Z(n831) );
  IVSVTX0H U986 ( .A(n748), .Z(n750) );
  F_ND2ASVTX2 U987 ( .A(n750), .B(n749), .Z(n829) );
  NR2SVTX0H U988 ( .A(n758), .B(n697), .Z(n759) );
  IVSVTX0H U989 ( .A(n765), .Z(n766) );
  AO7NSVTX1 U990 ( .A(n768), .B(n767), .C(n766), .Z(n769) );
  EOSVTX0H U991 ( .A(n770), .B(n769), .Z(n772) );
  NR2SVTX2 U992 ( .A(n774), .B(n773), .Z(n818) );
  FA1SVTX4 U993 ( .A(n780), .B(n779), .CI(n778), .CO(n785), .Z(n781) );
  IVSVTX2 U994 ( .A(n908), .Z(n783) );
  FA1SVTX1 U995 ( .A(n791), .B(n790), .CI(n789), .CO(n796), .Z(n792) );
  IVSVTX2 U996 ( .A(n815), .Z(n794) );
  IVSVTX0H U997 ( .A(n803), .Z(n806) );
  F_EOSVTX2 U998 ( .A(n804), .B(n915), .Z(O[25]) );
  IVSVTX0H U999 ( .A(n809), .Z(n810) );
  ND2SVTX2 U1000 ( .A(n811), .B(n810), .Z(n813) );
  F_EOSVTX2 U1001 ( .A(n813), .B(n812), .Z(O[23]) );
  IVSVTX0H U1002 ( .A(n818), .Z(n819) );
  IVSVTX0H U1003 ( .A(n823), .Z(n824) );
  IVSVTX0H U1004 ( .A(n832), .Z(n833) );
  IVSVTX0H U1005 ( .A(n837), .Z(n838) );
  IVSVTX0H U1006 ( .A(n841), .Z(n844) );
  IVSVTX0H U1007 ( .A(n842), .Z(n843) );
  AO6SVTX1 U1008 ( .A(n860), .B(n844), .C(n843), .Z(n845) );
  AO6SVTX1 U1009 ( .A(n860), .B(n850), .C(n849), .Z(n851) );
  IVSVTX0H U1010 ( .A(n862), .Z(n863) );
  AO7SVTX1 U1011 ( .A(n871), .B(n886), .C(n870), .Z(n882) );
  AO6SVTX1 U1012 ( .A(n882), .B(n880), .C(n872), .Z(n873) );
  AO7SVTX1 U1013 ( .A(n877), .B(n886), .C(n885), .Z(n878) );
  IVSVTX0H U1014 ( .A(n892), .Z(n893) );
  IVSVTX0H U1015 ( .A(n895), .Z(n901) );
  AO7SVTX1 U1016 ( .A(n898), .B(n901), .C(n900), .Z(n896) );
  IVSVTX0H U1017 ( .A(n898), .Z(n899) );
  IVSVTX0H U1018 ( .A(n903), .Z(n904) );
  AO7SVTX1 U1019 ( .A(n912), .B(n211), .C(n911), .Z(n914) );
endmodule

