
module m_rangemapping ( N, O );
  input [31:0] N;
  output [31:0] O;
  wire   n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n421, n422, n423, n424,
         n425, n426, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1763;

  BFSVTX0H U296 ( .A(n1221), .Z(O[28]) );
  IVSVTX0H U297 ( .A(n1569), .Z(n913) );
  IVSVTX0H U298 ( .A(n1626), .Z(n1629) );
  B_ND2SVTX2 U299 ( .A(n915), .B(n451), .Z(n1630) );
  F_ND2SVTX0H U300 ( .A(n1697), .B(n412), .Z(n1733) );
  B_ND2SVTX0H U301 ( .A(n1745), .B(n443), .Z(n1746) );
  BFSVTX4 U302 ( .A(n1614), .Z(n1616) );
  IVSVTX0H U303 ( .A(n1726), .Z(n1727) );
  IVSVTX2 U304 ( .A(n1621), .Z(n915) );
  IVSVTX0H U305 ( .A(n1711), .Z(n1713) );
  IVSVTX0H U306 ( .A(n790), .Z(n1756) );
  IVSVTX0H U307 ( .A(n1745), .Z(n1741) );
  IVSVTX0H U308 ( .A(n404), .Z(n1748) );
  IVSVTX0H U309 ( .A(n1687), .Z(n880) );
  IVSVTX0H U310 ( .A(n246), .Z(n907) );
  BFSVTX0H U311 ( .A(n1731), .Z(n412) );
  IVSVTX2 U312 ( .A(n1620), .Z(n451) );
  IVSVTX0H U313 ( .A(n462), .Z(n1712) );
  IVSVTX0H U314 ( .A(n1550), .Z(n528) );
  IVSVTX2 U315 ( .A(n937), .Z(n246) );
  IVSVTX0H U316 ( .A(n1674), .Z(n902) );
  BFSVTX0H U317 ( .A(n687), .Z(n686) );
  BFSVTX0H U318 ( .A(n1688), .Z(n436) );
  BFSVTX0H U319 ( .A(n1703), .Z(n462) );
  BFSVTX0H U320 ( .A(n1709), .Z(n483) );
  BFSVTX4 U321 ( .A(n1605), .Z(n1612) );
  BFSVTX0H U322 ( .A(n1652), .Z(n327) );
  BFSVTX2 U323 ( .A(n1702), .Z(n1710) );
  OR2SVTX2 U324 ( .A(n1496), .B(n1495), .Z(n937) );
  BFSVTX2 U325 ( .A(n1664), .Z(n1677) );
  NR2SVTX4 U326 ( .A(n926), .B(n1596), .Z(n1605) );
  ND2SVTX6 U327 ( .A(n1595), .B(n1594), .Z(n624) );
  IVSVTX2 U328 ( .A(n1514), .Z(n1593) );
  IVSVTX1 U329 ( .A(n229), .Z(n627) );
  CTIVSVTX2 U330 ( .A(n1586), .Z(n881) );
  ENSVTX1 U331 ( .A(n1498), .B(n1497), .Z(n736) );
  ND2SVTX6 U332 ( .A(n1503), .B(n738), .Z(n575) );
  AO5NSVTX4 U333 ( .A(n1572), .B(n1570), .C(n1571), .Z(n930) );
  AO4SVTX4 U334 ( .A(n1566), .B(n592), .C(n920), .D(n633), .Z(n591) );
  IVSVTX2 U335 ( .A(n771), .Z(n1570) );
  B_IVSVTX1 U336 ( .A(n883), .Z(n939) );
  F_ENSVTX2 U337 ( .A(n457), .B(n230), .Z(n1526) );
  IVSVTX2 U338 ( .A(n604), .Z(n631) );
  ND3SVTX6 U339 ( .A(n1513), .B(n1512), .C(n1511), .Z(n1585) );
  NR3SVTX4 U340 ( .A(n496), .B(n1578), .C(n873), .Z(n580) );
  ENSVTX0H U341 ( .A(n770), .B(n877), .Z(n772) );
  ENSVTX2 U342 ( .A(n651), .B(n1500), .Z(n1505) );
  IVSVTX0H U343 ( .A(n445), .Z(n1556) );
  AO2ABSVTX6 U344 ( .C(n873), .D(n623), .A(n249), .B(n1576), .Z(n452) );
  ENSVTX0H U345 ( .A(n648), .B(n1499), .Z(n651) );
  HA1SVTX1 U346 ( .A(n322), .B(n1545), .CO(n1575), .S(n1572) );
  IVSVTX0H U347 ( .A(n1528), .Z(n1530) );
  IVSVTX2 U348 ( .A(n876), .Z(n877) );
  IVSVTX0H U349 ( .A(n922), .Z(n470) );
  FAS1SVTX2 U350 ( .A(n1245), .B(n1502), .CI(n1501), .CO(n1500), .Z(n1527) );
  IVSVTX10 U351 ( .A(n1578), .Z(n1521) );
  IVSVTX0H U352 ( .A(n1546), .Z(n1547) );
  IVSVTX0H U353 ( .A(n1554), .Z(n876) );
  BFSVTX2 U354 ( .A(n1660), .Z(n1553) );
  IVSVTX0H U355 ( .A(n1507), .Z(n1306) );
  F_AN2SVTX2 U356 ( .A(n448), .B(n684), .Z(n1546) );
  BFSVTX2 U357 ( .A(n1529), .Z(n447) );
  IVSVTX0H U358 ( .A(n1532), .Z(n1557) );
  BFSVTX2 U359 ( .A(n1558), .Z(n449) );
  BFSVTX0H U360 ( .A(n417), .Z(n448) );
  IVSVTX0H U361 ( .A(n1549), .Z(n1661) );
  ND2SVTX2 U362 ( .A(n1498), .B(n1491), .Z(n620) );
  F_ND2SVTX1 U363 ( .A(n1498), .B(n1490), .Z(n618) );
  NR2SVTX4 U364 ( .A(n1507), .B(n1582), .Z(n1490) );
  BFSVTX2 U365 ( .A(n1533), .Z(n1559) );
  NR2SVTX6 U366 ( .A(n1507), .B(n1581), .Z(n1491) );
  NR2SVTX6 U367 ( .A(n1532), .B(n539), .Z(n1508) );
  NR2ASVTX6 U368 ( .A(n603), .B(n1499), .Z(n1507) );
  AO6SVTX6 U369 ( .A(n1551), .B(n1308), .C(n1292), .Z(n1536) );
  NR2ASVTX4 U370 ( .A(n289), .B(n1501), .Z(n1581) );
  IVSVTX2 U371 ( .A(n220), .Z(n247) );
  CTIVSVTX2 U372 ( .A(n1291), .Z(n782) );
  NR2SVTX6 U373 ( .A(n1534), .B(n1528), .Z(n845) );
  AO3SVTX6 U374 ( .A(n1474), .B(n1703), .C(n1473), .D(n1701), .Z(n1667) );
  ND2SVTX4 U375 ( .A(n1758), .B(n1421), .Z(n1423) );
  ND2SVTX6 U376 ( .A(n919), .B(n1664), .Z(n1484) );
  ND2ASVTX6 U377 ( .A(n1451), .B(n279), .Z(n1716) );
  ND2ASVTX6 U378 ( .A(n460), .B(n1358), .Z(n1652) );
  BFSVTX6 U379 ( .A(n1686), .Z(n461) );
  IVSVTX0H U380 ( .A(n253), .Z(n1294) );
  IVSVTX4 U381 ( .A(n1454), .Z(n281) );
  IVSVTX4 U382 ( .A(n1672), .Z(n1482) );
  IVSVTX2 U383 ( .A(n1447), .Z(n670) );
  ND2ASVTX6 U384 ( .A(n236), .B(n841), .Z(n1688) );
  NR2SVTX2 U385 ( .A(n547), .B(n1409), .Z(n546) );
  IVSVTX4 U386 ( .A(n410), .Z(n1383) );
  IVSVTX4 U387 ( .A(n1686), .Z(n1478) );
  AO2ABSVTX6 U388 ( .C(n586), .D(n698), .A(n654), .B(n875), .Z(n587) );
  IVSVTX4 U389 ( .A(n763), .Z(n761) );
  AO2SVTX4 U390 ( .A(n767), .B(n921), .C(n840), .D(n849), .Z(n848) );
  AO2ABSVTX6 U391 ( .C(n921), .D(n1246), .A(n875), .B(n230), .Z(n809) );
  ND2SVTX4 U392 ( .A(n874), .B(n1288), .Z(n798) );
  ND2ASVTX6 U393 ( .A(n1285), .B(n740), .Z(n704) );
  ND2ASVTX6 U394 ( .A(n1476), .B(n726), .Z(n455) );
  IVSVTX0H U395 ( .A(n754), .Z(n1399) );
  IVSVTX2 U396 ( .A(n251), .Z(n840) );
  IVSVTX2 U397 ( .A(n478), .Z(n331) );
  IVSVTX0H U398 ( .A(n1467), .Z(n316) );
  ND2ASVTX4 U399 ( .A(n289), .B(n741), .Z(n601) );
  IVSVTX0H U400 ( .A(n1419), .Z(n256) );
  IVSVTX12 U401 ( .A(n836), .Z(n873) );
  IVSVTX2 U402 ( .A(n856), .Z(n252) );
  IVSVTX2 U403 ( .A(n887), .Z(n1406) );
  ND2ASVTX6 U404 ( .A(n478), .B(n1352), .Z(n1460) );
  ND2ASVTX6 U405 ( .A(n1443), .B(n1376), .Z(n1477) );
  IVSVTX2 U406 ( .A(n1285), .Z(n802) );
  IVSVTX2 U407 ( .A(n1410), .Z(n889) );
  ND2ASVTX6 U408 ( .A(n1443), .B(n1322), .Z(n751) );
  IVSVTX4 U409 ( .A(n1577), .Z(n1353) );
  IVSVTX4 U410 ( .A(n1515), .Z(n230) );
  IVSVTX2 U411 ( .A(n1438), .Z(n1439) );
  CTIVSVTX2 U412 ( .A(n652), .Z(n1428) );
  AO6SVTX4 U413 ( .A(n1441), .B(n874), .C(n1440), .Z(n1445) );
  BFSVTX6 U414 ( .A(n1498), .Z(n675) );
  NR2ASVTX4 U415 ( .A(n1480), .B(n875), .Z(n1476) );
  ND2ASVTX4 U416 ( .A(n1248), .B(n225), .Z(n750) );
  IVSVTX0H U417 ( .A(n238), .Z(n1467) );
  IVSVTX4 U418 ( .A(n232), .Z(n884) );
  ND2SVTX6 U419 ( .A(n770), .B(n213), .Z(n707) );
  ND2SVTX4 U420 ( .A(n645), .B(n1403), .Z(n374) );
  IVSVTX4 U421 ( .A(n740), .Z(n701) );
  IVSVTX6 U422 ( .A(n855), .Z(n640) );
  BFSVTX4 U423 ( .A(n1436), .Z(n478) );
  IVSVTX6 U424 ( .A(n1248), .Z(n232) );
  NR2SVTX2 U425 ( .A(n237), .B(n534), .Z(n1321) );
  CTIVSVTX2 U426 ( .A(n584), .Z(n560) );
  IVSVTX2 U427 ( .A(n1466), .Z(n238) );
  NR2SVTX2 U428 ( .A(n1420), .B(n521), .Z(n844) );
  IVSVTX4 U429 ( .A(n832), .Z(n1380) );
  NR2SVTX4 U430 ( .A(n684), .B(n417), .Z(n378) );
  AO7SVTX4 U431 ( .A(n1245), .B(n743), .C(n1299), .Z(n1239) );
  EOSVTX4 U432 ( .A(n754), .B(n1433), .Z(n1403) );
  NR2ASVTX4 U433 ( .A(n1373), .B(n875), .Z(n1374) );
  IVSVTX8 U434 ( .A(n534), .Z(n249) );
  CTBUFSVTX4 U435 ( .A(n1436), .Z(n521) );
  IVSVTX8 U436 ( .A(n654), .Z(n1519) );
  IVSVTX2 U437 ( .A(n1047), .Z(n1510) );
  IVSVTX10 U438 ( .A(n578), .Z(n875) );
  IVSVTX2 U439 ( .A(n1299), .Z(n603) );
  IVSVTX10 U440 ( .A(n1577), .Z(n1443) );
  IVSVTX2 U441 ( .A(n1451), .Z(n1453) );
  IVSVTX8 U442 ( .A(n684), .Z(n920) );
  IVSVTX0H U443 ( .A(n1386), .Z(n1387) );
  IVSVTX1 U444 ( .A(n424), .Z(n1045) );
  F_IVSVTX1 U445 ( .A(n1461), .Z(n1427) );
  NR2SVTX6 U446 ( .A(n754), .B(n1433), .Z(n787) );
  ND2ASVTX4 U447 ( .A(n1339), .B(n1330), .Z(n1475) );
  IVSVTX8 U448 ( .A(n872), .Z(n836) );
  IVSVTX2 U449 ( .A(n1420), .Z(n403) );
  F_ND2ASVTX2 U450 ( .A(n497), .B(n1182), .Z(n1466) );
  CTIVSVTX6 U451 ( .A(n1289), .Z(n251) );
  IVSVTX2 U452 ( .A(n1458), .Z(n1429) );
  CTBUFSVTX4 U453 ( .A(n1424), .Z(n468) );
  BFSVTX0H U454 ( .A(n1384), .Z(n317) );
  BFSVTX8 U455 ( .A(n1230), .Z(n684) );
  IVSVTX2 U456 ( .A(n418), .Z(n1425) );
  IVSVTX2 U457 ( .A(n1349), .Z(n1330) );
  IVSVTX2 U458 ( .A(n1360), .Z(n569) );
  IVSVTX10 U459 ( .A(n1433), .Z(n1398) );
  NR2SVTX6 U460 ( .A(n866), .B(n1229), .Z(n605) );
  NR2SVTX4 U461 ( .A(n1141), .B(n362), .Z(n348) );
  IVSVTX6 U462 ( .A(n1245), .Z(n289) );
  IVSVTX8 U463 ( .A(n1436), .Z(n1577) );
  ND2SVTX1 U464 ( .A(n729), .B(n274), .Z(n932) );
  NR2SVTX2 U465 ( .A(n424), .B(n1273), .Z(n490) );
  B_IVSVTX1 U466 ( .A(n500), .Z(n582) );
  CTIVSVTX6 U467 ( .A(n1373), .Z(n306) );
  IVSVTX2 U468 ( .A(n1424), .Z(n491) );
  IVSVTX2 U469 ( .A(n1311), .Z(n1336) );
  ND2SVTX2 U470 ( .A(n1182), .B(n825), .Z(n1337) );
  AO7SVTX4 U471 ( .A(n424), .B(n1323), .C(n1319), .Z(n1468) );
  ND3ASVTX4 U472 ( .A(n1338), .B(n1348), .C(n1426), .Z(n492) );
  ND2SVTX4 U473 ( .A(n1251), .B(n1235), .Z(n804) );
  NR2SVTX6 U474 ( .A(n1480), .B(n1360), .Z(n555) );
  F_ND2ASVTX2 U475 ( .A(n294), .B(n274), .Z(n898) );
  IVSVTX0H U476 ( .A(n1389), .Z(n1391) );
  NR2ASVTX1 U477 ( .A(n1388), .B(n233), .Z(n1392) );
  AN2SVTX6 U478 ( .A(n803), .B(n1074), .Z(n925) );
  ND2SVTX4 U479 ( .A(n766), .B(n510), .Z(n507) );
  IVSVTX2 U480 ( .A(n1361), .Z(n764) );
  NR3SVTX4 U481 ( .A(n350), .B(n1390), .C(n1281), .Z(n1284) );
  ND2ASVTX4 U482 ( .A(n885), .B(n826), .Z(n1096) );
  NR2SVTX2 U483 ( .A(n1184), .B(n1185), .Z(n1075) );
  IVSVTX4 U484 ( .A(n1232), .Z(n671) );
  CTBUFSVTX4 U485 ( .A(n1397), .Z(n431) );
  BFSVTX8 U486 ( .A(n1390), .Z(n424) );
  NR2ASVTX6 U487 ( .A(n1277), .B(n765), .Z(n1362) );
  IVSVTX2 U488 ( .A(n1181), .Z(n810) );
  B_IVSVTX1 U489 ( .A(n1346), .Z(n211) );
  AN3BCSVTX4 U490 ( .A(n1251), .B(n904), .C(n1052), .Z(n1361) );
  ND2SVTX6 U491 ( .A(n1093), .B(n239), .Z(n635) );
  ND4ABSVTX6 U492 ( .A(n1211), .B(n1212), .C(n1210), .D(n1209), .Z(n425) );
  IVSVTX4 U493 ( .A(n341), .Z(n497) );
  IVSVTX4 U494 ( .A(n362), .Z(n356) );
  AO4SVTX4 U495 ( .A(n302), .B(n1184), .C(n1108), .D(n1109), .Z(n275) );
  AO6ASVTX6 U496 ( .A(n933), .B(n297), .C(n222), .Z(n1080) );
  AO4SVTX6 U497 ( .A(n1183), .B(n1184), .C(n1109), .D(n1185), .Z(n509) );
  ND2ASVTX4 U498 ( .A(n241), .B(n1236), .Z(n1110) );
  IVSVTX2 U499 ( .A(n231), .Z(n480) );
  BFSVTX4 U500 ( .A(n1107), .Z(n302) );
  F_IVSVTX1 U501 ( .A(n387), .Z(n933) );
  IVSVTX2 U502 ( .A(n1094), .Z(n1185) );
  ND2SVTX2 U503 ( .A(n778), .B(n830), .Z(n471) );
  ND3SVTX6 U504 ( .A(n1043), .B(n1044), .C(n685), .Z(n673) );
  CTIVSVTX6 U505 ( .A(n1273), .Z(n329) );
  ND2SVTX4 U506 ( .A(n885), .B(n1261), .Z(n341) );
  AO7SVTX6 U507 ( .A(n838), .B(n435), .C(n837), .Z(n285) );
  IVSVTX4 U508 ( .A(n269), .Z(n1407) );
  ND4ABSVTX4 U509 ( .A(n1211), .B(n1212), .C(n1210), .D(n1209), .Z(n1260) );
  CTIVSVTX2 U510 ( .A(n1163), .Z(n1167) );
  NR2SVTX2 U511 ( .A(n1103), .B(n1184), .Z(n1106) );
  IVSVTX4 U512 ( .A(n1390), .Z(O[27]) );
  NR2SVTX4 U513 ( .A(n1251), .B(n1042), .Z(n685) );
  ND2SVTX2 U514 ( .A(n1056), .B(n1057), .Z(n1077) );
  ND2SVTX6 U515 ( .A(n690), .B(n1040), .Z(n1093) );
  ND3ABSVTX6 U516 ( .A(n747), .B(n242), .C(n1221), .Z(n1327) );
  ND2SVTX4 U517 ( .A(n1130), .B(n1397), .Z(n1128) );
  AO2SVTX4 U518 ( .A(n274), .B(n1099), .C(n240), .D(n1100), .Z(n1101) );
  CTIVSVTX2 U519 ( .A(n778), .Z(n1183) );
  BFSVTX6 U520 ( .A(n371), .Z(n435) );
  BFSVTX6 U521 ( .A(n1411), .Z(n428) );
  NR2ASVTX6 U522 ( .A(n545), .B(n1132), .Z(n296) );
  NR2SVTX2 U523 ( .A(n815), .B(n1215), .Z(n381) );
  IVSVTX8 U524 ( .A(n885), .Z(n766) );
  IVSVTX2 U525 ( .A(n1042), .Z(n543) );
  ND3SVTX4 U526 ( .A(n1254), .B(n226), .C(n1192), .Z(n514) );
  NR2ASVTX4 U527 ( .A(n815), .B(n1223), .Z(n551) );
  ND2ASVTX4 U528 ( .A(n1162), .B(n1203), .Z(n1316) );
  AO7SVTX1 U529 ( .A(n961), .B(n1069), .C(n235), .Z(n962) );
  ND3SVTX4 U530 ( .A(n1334), .B(n485), .C(n1333), .Z(n611) );
  BFSVTX4 U531 ( .A(n904), .Z(n326) );
  IVSVTX10 U532 ( .A(n486), .Z(n1109) );
  CTIVSVTX2 U533 ( .A(n1180), .Z(n1168) );
  IVSVTX2 U534 ( .A(n664), .Z(n662) );
  IVSVTX0H U535 ( .A(n259), .Z(n734) );
  ND2SVTX4 U536 ( .A(n1033), .B(n1032), .Z(n1100) );
  IVSVTX8 U537 ( .A(n1411), .Z(n885) );
  ND3SVTX4 U538 ( .A(n717), .B(n1214), .C(n233), .Z(n711) );
  CTIVSVTX2 U539 ( .A(n1402), .Z(n733) );
  AO6SVTX2 U540 ( .A(n1196), .B(n815), .C(n1174), .Z(n1148) );
  ND3SVTX6 U541 ( .A(n1048), .B(n1049), .C(n792), .Z(n1037) );
  AO6SVTX6 U542 ( .A(n683), .B(n1188), .C(n1055), .Z(n777) );
  ND3SVTX4 U543 ( .A(n1267), .B(n714), .C(n545), .Z(n713) );
  AO6ASVTX2 U544 ( .A(n1058), .B(n595), .C(n916), .Z(n661) );
  IVSVTX2 U545 ( .A(n1206), .Z(n1325) );
  BFSVTX10 U546 ( .A(n385), .Z(n350) );
  BFSVTX10 U547 ( .A(n892), .Z(n1390) );
  IVSVTX2 U548 ( .A(n897), .Z(n865) );
  NR2SVTX2 U549 ( .A(n1280), .B(n924), .Z(n863) );
  IVSVTX0H U550 ( .A(n262), .Z(n1129) );
  AN3SVTX4 U551 ( .A(n1034), .B(n815), .C(n957), .Z(n935) );
  NR2ASVTX4 U552 ( .A(n1178), .B(n786), .Z(n664) );
  AO6ABSVTX6 U553 ( .A(n941), .B(n682), .C(n1177), .Z(n1204) );
  AO7ASVTX2 U554 ( .A(N[12]), .B(n959), .C(n1002), .Z(n916) );
  NR2SVTX2 U555 ( .A(n965), .B(n964), .Z(n966) );
  ND2SVTX2 U556 ( .A(n1144), .B(n1169), .Z(n1170) );
  ND3ASVTX4 U557 ( .A(n1118), .B(n258), .C(n1036), .Z(n1048) );
  ND2SVTX6 U558 ( .A(n1063), .B(n1062), .Z(n1094) );
  AO6ASVTX4 U559 ( .A(n958), .B(n663), .C(n1003), .Z(n1056) );
  ND2ASVTX4 U560 ( .A(n262), .B(n1004), .Z(n967) );
  CTIVSVTX2 U561 ( .A(n242), .Z(n345) );
  ND3ABSVTX4 U562 ( .A(n1172), .B(n1118), .C(n293), .Z(n1119) );
  IVSVTX12 U563 ( .A(n1041), .Z(n1205) );
  F_ND2ASVTX2 U564 ( .A(n775), .B(n663), .Z(n1032) );
  IVSVTX2 U565 ( .A(n959), .Z(n1036) );
  AO6SVTX1 U566 ( .A(n776), .B(N[1]), .C(n1068), .Z(n775) );
  AO7SVTX4 U567 ( .A(n1195), .B(n853), .C(n1280), .Z(n1206) );
  ND2ASVTX6 U568 ( .A(n1171), .B(n1144), .Z(n1196) );
  IVSVTX2 U569 ( .A(n1177), .Z(n1202) );
  IVSVTX6 U570 ( .A(n266), .Z(n540) );
  F_AO7ASVTX1 U571 ( .A(n1151), .B(n959), .C(n1030), .Z(n1031) );
  IVSVTX6 U572 ( .A(n691), .Z(n1186) );
  IVSVTX10 U573 ( .A(n999), .Z(n683) );
  IVSVTX2 U574 ( .A(n383), .Z(n382) );
  IVSVTX2 U575 ( .A(n1125), .Z(n897) );
  IVSVTX2 U576 ( .A(n1136), .Z(n259) );
  IVSVTX2 U577 ( .A(n257), .Z(n882) );
  NR2ASVTX4 U578 ( .A(n827), .B(n1160), .Z(n1215) );
  IVSVTX0H U579 ( .A(N[7]), .Z(n1118) );
  CTIVSVTX4 U580 ( .A(n1280), .Z(O[29]) );
  IVSVTX4 U581 ( .A(n1314), .Z(n1223) );
  IVSVTX0H U582 ( .A(n245), .Z(n829) );
  ND2ASVTX4 U583 ( .A(n1389), .B(n358), .Z(n402) );
  IVSVTX4 U584 ( .A(n892), .Z(n415) );
  NR2ASVTX2 U585 ( .A(N[18]), .B(n258), .Z(n965) );
  NR2SVTX2 U586 ( .A(n1146), .B(n1172), .Z(n409) );
  AO6CSVTX6 U587 ( .A(n595), .B(n594), .C(n1073), .Z(n716) );
  NR2ASVTX2 U588 ( .A(n918), .B(n1059), .Z(n1063) );
  ND2SVTX1 U589 ( .A(n245), .B(n776), .Z(n1034) );
  ND2SVTX1 U590 ( .A(N[2]), .B(n1145), .Z(n749) );
  ND2ASVTX6 U591 ( .A(n272), .B(n731), .Z(n271) );
  NR2ASVTX4 U592 ( .A(n594), .B(n1172), .Z(n1171) );
  AN3SVTX6 U593 ( .A(n386), .B(N[12]), .C(n258), .Z(n1177) );
  IVSVTX2 U594 ( .A(n827), .Z(n1161) );
  BFSVTX0H U595 ( .A(n1000), .Z(n1001) );
  AN3CSVTX4 U596 ( .A(n1150), .B(n337), .C(n824), .Z(n1180) );
  ND3ABSVTX4 U597 ( .A(n262), .B(n493), .C(n1084), .Z(n1144) );
  NR3SVTX4 U598 ( .A(n262), .B(n959), .C(n960), .Z(n718) );
  ND2ASVTX4 U599 ( .A(N[2]), .B(n1134), .Z(n753) );
  NR2ASVTX2 U600 ( .A(n1178), .B(n1069), .Z(n1059) );
  IVSVTX4 U601 ( .A(n293), .Z(n361) );
  CTIVSVTX2 U602 ( .A(n298), .Z(n896) );
  IVSVTX2 U603 ( .A(n1116), .Z(n552) );
  ND2SVTX2 U604 ( .A(n989), .B(n493), .Z(n494) );
  IVSVTX0H U605 ( .A(n261), .Z(n272) );
  F_ND2ASVTX2 U606 ( .A(n1146), .B(n1145), .Z(n822) );
  ND2SVTX2 U607 ( .A(n258), .B(n1086), .Z(n1090) );
  F_ND2SVTX1 U608 ( .A(n235), .B(n800), .Z(n824) );
  ND2SVTX2 U609 ( .A(n1188), .B(n493), .Z(n1216) );
  IVSVTX0H U610 ( .A(n1068), .Z(n517) );
  B_ND2SVTX2 U611 ( .A(N[4]), .B(n1154), .Z(n1124) );
  IVSVTX4 U612 ( .A(n1172), .Z(n666) );
  ND2SVTX2 U613 ( .A(N[0]), .B(n1145), .Z(n1123) );
  BFSVTX0H U614 ( .A(N[4]), .Z(n1178) );
  NR2ASVTX2 U615 ( .A(N[5]), .B(n776), .Z(n1189) );
  BFSVTX4 U616 ( .A(n1143), .Z(n493) );
  IVSVTX0H U617 ( .A(n958), .Z(n1088) );
  ND2ASVTX6 U618 ( .A(n261), .B(n1172), .Z(n1152) );
  ND2SVTX2 U619 ( .A(n1021), .B(n235), .Z(n1022) );
  F_IVSVTX1 U620 ( .A(n1016), .Z(n1017) );
  IVSVTX2 U621 ( .A(N[1]), .Z(n261) );
  ND2SVTX4 U622 ( .A(n821), .B(n818), .Z(n816) );
  IVSVTX2 U623 ( .A(n820), .Z(n817) );
  ND3SVTX4 U624 ( .A(n393), .B(n392), .C(n391), .Z(n390) );
  IVSVTX6 U625 ( .A(n912), .Z(n1153) );
  IVSVTX2 U626 ( .A(n894), .Z(n235) );
  NR4SVTX4 U627 ( .A(n667), .B(n956), .C(n955), .D(n446), .Z(n818) );
  NR3SVTX4 U628 ( .A(n1135), .B(n992), .C(n991), .Z(n392) );
  ND2SVTX2 U629 ( .A(n1026), .B(n1068), .Z(n1027) );
  AO7SVTX2 U630 ( .A(n422), .B(n970), .C(n398), .Z(n397) );
  IVSVTX2 U631 ( .A(n947), .Z(n986) );
  F_IVSVTX1 U632 ( .A(n945), .Z(n894) );
  BFSVTX4 U633 ( .A(n1023), .Z(n437) );
  NR3SVTX4 U634 ( .A(n1085), .B(N[7]), .C(n990), .Z(n944) );
  AO6SVTX4 U635 ( .A(n1010), .B(n594), .C(n989), .Z(n995) );
  IVSVTX6 U636 ( .A(N[27]), .Z(n957) );
  NR2ASVTX2 U637 ( .A(N[18]), .B(n422), .Z(n988) );
  IVSVTX2 U638 ( .A(n992), .Z(n793) );
  ND2ASVTX6 U639 ( .A(N[29]), .B(n851), .Z(n972) );
  IVSVTX4 U640 ( .A(n943), .Z(n1010) );
  IVSVTX4 U641 ( .A(n989), .Z(n961) );
  IVSVTX4 U642 ( .A(N[22]), .Z(n1039) );
  ND2ASVTX6 U643 ( .A(N[8]), .B(n263), .Z(n949) );
  ND2SVTX2 U644 ( .A(n369), .B(n475), .Z(n975) );
  BFSVTX4 U645 ( .A(N[29]), .Z(n1021) );
  CTBUFSVTX4 U646 ( .A(N[28]), .Z(n1000) );
  IVSVTX4 U647 ( .A(n973), .Z(n991) );
  IVSVTX4 U648 ( .A(N[2]), .Z(n262) );
  IVSVTX4 U649 ( .A(N[6]), .Z(n1146) );
  ND2SVTX4 U650 ( .A(n1005), .B(n1008), .Z(n979) );
  NR2SVTX6 U651 ( .A(N[27]), .B(N[24]), .Z(n769) );
  IVSVTX8 U652 ( .A(N[24]), .Z(n475) );
  NR2SVTX6 U653 ( .A(N[19]), .B(N[29]), .Z(n369) );
  NR2SVTX6 U654 ( .A(N[17]), .B(N[16]), .Z(n368) );
  IVSVTX4 U655 ( .A(N[13]), .Z(n1005) );
  NR2SVTX4 U656 ( .A(N[27]), .B(N[25]), .Z(n346) );
  CTIVSVTX6 U657 ( .A(n511), .Z(n1576) );
  MUX21NSVTX6 U658 ( .A(n922), .B(n911), .S(n1576), .Z(n1580) );
  ND3ABSVTX8 U659 ( .A(n1300), .B(n675), .C(n681), .Z(n680) );
  ENSVTX8 U660 ( .A(n1377), .B(n487), .Z(n1355) );
  NR4ABSVTX6 U661 ( .A(n309), .B(n1345), .C(n211), .D(n1344), .Z(n1347) );
  AO7SVTX4 U662 ( .A(n677), .B(n678), .C(n1241), .Z(n1242) );
  ND3SVTX6 U663 ( .A(n212), .B(n1066), .C(n1065), .Z(n1235) );
  ND2SVTX4 U664 ( .A(n1094), .B(n891), .Z(n212) );
  ND2ASVTX8 U665 ( .A(n770), .B(n640), .Z(n858) );
  IVSVTX12 U666 ( .A(n724), .Z(n266) );
  AO6SVTX4 U667 ( .A(n1578), .B(n470), .C(n911), .Z(n1511) );
  BFSVTX4 U668 ( .A(n1293), .Z(n213) );
  NR2SVTX6 U669 ( .A(n1618), .B(n1620), .Z(n1614) );
  F_IVSVTX1 U670 ( .A(n1581), .Z(n334) );
  F_IVSVTX1 U671 ( .A(n1353), .Z(n911) );
  AO3ABSVTX6 U672 ( .A(n1299), .B(n695), .C(n1239), .D(n873), .Z(n677) );
  AO7ABSVTX6 U673 ( .A(n921), .B(n225), .C(n1432), .Z(n1452) );
  ND3SVTX6 U674 ( .A(n1426), .B(n1425), .C(n468), .Z(n854) );
  ND2SVTX6 U675 ( .A(n993), .B(n1016), .Z(n994) );
  NR2SVTX6 U676 ( .A(n1401), .B(n294), .Z(n295) );
  ND2ASVTX8 U677 ( .A(n1245), .B(n763), .Z(n762) );
  ND2ASVTX8 U678 ( .A(n723), .B(n1271), .Z(n1289) );
  IVSVTX8 U679 ( .A(n511), .Z(n495) );
  IVSVTX12 U680 ( .A(n495), .Z(n496) );
  AO7SVTX8 U681 ( .A(n1660), .B(n1291), .C(n1290), .Z(n1292) );
  ENSVTX4 U682 ( .A(n736), .B(n575), .Z(n1597) );
  ENSVTX8 U683 ( .A(n1429), .B(n481), .Z(n1435) );
  BFSVTX6 U684 ( .A(n1695), .Z(n214) );
  ENSVTX6 U685 ( .A(n567), .B(n571), .Z(n1359) );
  IVSVTX4 U686 ( .A(n215), .Z(n227) );
  ND2SVTX4 U687 ( .A(n699), .B(n286), .Z(n215) );
  AO6CSVTX2 U688 ( .A(N[1]), .B(n776), .C(n517), .Z(n518) );
  IVSVTX0H U689 ( .A(n1137), .Z(n553) );
  NR2SVTX2 U690 ( .A(n289), .B(n695), .Z(n1243) );
  ND2SVTX2 U691 ( .A(N[5]), .B(n1153), .Z(n360) );
  AO7NSVTX4 U692 ( .A(n1087), .B(n682), .C(n1089), .Z(n934) );
  NR2SVTX2 U693 ( .A(n1146), .B(n786), .Z(n963) );
  IVSVTX0H U694 ( .A(n1198), .Z(n1162) );
  AO2SVTX6 U695 ( .A(n545), .B(n515), .C(n1203), .D(n221), .Z(n1192) );
  ND2SVTX2 U696 ( .A(n830), .B(n1077), .Z(n1079) );
  IVSVTX2 U697 ( .A(n1165), .Z(n1166) );
  AO7SVTX6 U698 ( .A(n1226), .B(n1225), .C(n799), .Z(n1346) );
  NR3SVTX6 U699 ( .A(n1047), .B(n1404), .C(n920), .Z(n377) );
  IVSVTX2 U700 ( .A(n1417), .Z(n254) );
  IVSVTX2 U701 ( .A(n635), .Z(n888) );
  IVSVTX0H U702 ( .A(n1306), .Z(n905) );
  IVSVTX0H U703 ( .A(n1697), .Z(n1730) );
  AO7SVTX4 U704 ( .A(n1612), .B(n1608), .C(n1607), .Z(n1609) );
  AO6SVTX1 U705 ( .A(n1759), .B(n1758), .C(n1757), .Z(n1760) );
  F_ND2SVTX0H U706 ( .A(n1728), .B(n1727), .Z(n1729) );
  EOSVTX1 U707 ( .A(n1746), .B(n923), .Z(O[2]) );
  AN3SVTX6 U708 ( .A(n920), .B(n417), .C(n707), .Z(n216) );
  AN2SVTX4 U709 ( .A(n1406), .B(n843), .Z(n217) );
  AO7NSVTX4 U710 ( .A(n1053), .B(n1084), .C(n1054), .Z(n218) );
  AN2SVTX6 U711 ( .A(n553), .B(n1084), .Z(n219) );
  AO3NSVTX8 U712 ( .A(n318), .B(n1353), .C(n857), .D(n250), .Z(n220) );
  IVSVTX4 U713 ( .A(n422), .Z(n244) );
  IVSVTX2 U714 ( .A(n1214), .Z(n1103) );
  AO7NSVTX6 U715 ( .A(n1199), .B(n896), .C(n815), .Z(n221) );
  IVSVTX8 U716 ( .A(n1763), .Z(n1280) );
  IVSVTX12 U717 ( .A(n1763), .Z(n814) );
  IVSVTX12 U718 ( .A(n258), .Z(n960) );
  IVSVTX4 U719 ( .A(n917), .Z(n1038) );
  IVSVTX2 U720 ( .A(n1069), .Z(n243) );
  AN2SVTX4 U721 ( .A(n1100), .B(n830), .Z(n222) );
  ND3SVTX4 U722 ( .A(n1168), .B(n1179), .C(n358), .Z(n597) );
  AO7NSVTX2 U723 ( .A(n1251), .B(n1334), .C(n1333), .Z(n223) );
  IVSVTX2 U724 ( .A(n385), .Z(n859) );
  OR2SVTX4 U725 ( .A(n238), .B(n875), .Z(n224) );
  EOSVTX8 U726 ( .A(n1466), .B(n1313), .Z(n225) );
  AO7NSVTX4 U727 ( .A(n1191), .B(n1187), .C(n1278), .Z(n226) );
  NR2ASVTX2 U728 ( .A(n1574), .B(n875), .Z(n1287) );
  F_AN2SVTX2 U729 ( .A(n624), .B(n1619), .Z(n228) );
  F_EOSVTX2 U730 ( .A(n772), .B(n1565), .Z(n229) );
  IVSVTX6 U731 ( .A(n985), .Z(n389) );
  AN2SVTX6 U732 ( .A(n728), .B(n399), .Z(n1426) );
  IVSVTX8 U733 ( .A(n336), .Z(n860) );
  MUX21NSVTX6 U734 ( .A(n431), .B(n1130), .S(n435), .Z(n1449) );
  ND3ABSVTX6 U735 ( .A(n1546), .B(n496), .C(n623), .Z(n738) );
  IVSVTX8 U736 ( .A(n783), .Z(n1220) );
  AO5SVTX2 U737 ( .A(n1586), .B(n631), .C(n1585), .Z(n1514) );
  ND2ASVTX8 U738 ( .A(n1546), .B(n1548), .Z(n1571) );
  AO7SVTX8 U739 ( .A(n1537), .B(n1528), .C(n1529), .Z(n1298) );
  ND2SVTX2 U740 ( .A(n873), .B(n1382), .Z(n847) );
  ND3SVTX8 U741 ( .A(n961), .B(n951), .C(n950), .Z(n954) );
  IVSVTX12 U742 ( .A(n541), .Z(n724) );
  IVSVTX10 U743 ( .A(n408), .Z(n748) );
  AO6CSVTX8 U744 ( .A(n1202), .B(n927), .C(n815), .Z(n1226) );
  NR2ASVTX6 U745 ( .A(n1247), .B(n1545), .Z(n807) );
  AO7SVTX8 U746 ( .A(n1632), .B(n1639), .C(n1633), .Z(n1590) );
  AO5ASVTX8 U747 ( .B(n477), .A(n1527), .C(n590), .Z(n926) );
  IVSVTX4 U748 ( .A(n1635), .Z(n1642) );
  AO6SVTX4 U749 ( .A(n1615), .B(n1599), .C(n1598), .Z(n1600) );
  ND2SVTX4 U750 ( .A(n929), .B(n1597), .Z(n1604) );
  CTIVSVTX2 U751 ( .A(n737), .Z(n929) );
  NR2SVTX6 U752 ( .A(n580), .B(n579), .Z(n590) );
  B_ND2SVTX2 U753 ( .A(n1492), .B(n1513), .Z(n1623) );
  ND2SVTX2 U754 ( .A(n1557), .B(n1540), .Z(n1542) );
  CTIVSVTX2 U755 ( .A(n1559), .Z(n1535) );
  B_ND2SVTX2 U756 ( .A(n648), .B(n1500), .Z(n650) );
  F_ENSVTX2 U757 ( .A(n1738), .B(n1737), .Z(O[4]) );
  F_ENSVTX2 U758 ( .A(n1743), .B(n1742), .Z(O[3]) );
  B_ND2SVTX2 U759 ( .A(n1701), .B(n1700), .Z(n1708) );
  AO6SVTX6 U760 ( .A(n1421), .B(n1757), .C(n476), .Z(n1422) );
  AO2SVTX4 U761 ( .A(n232), .B(n1410), .C(n578), .D(n1419), .Z(n577) );
  IVSVTX10 U762 ( .A(n766), .Z(n231) );
  AO7SVTX4 U763 ( .A(n261), .B(n1159), .C(n1122), .Z(n1125) );
  AO7SVTX4 U764 ( .A(n1602), .B(n1607), .C(n1604), .Z(n1598) );
  B_ND2SVTX2 U765 ( .A(n1634), .B(n1633), .Z(n1637) );
  F_ND2ASVTX2 U766 ( .A(n229), .B(n1567), .Z(n1649) );
  NR2ASVTX2 U767 ( .A(n229), .B(n1567), .Z(n1647) );
  ND2SVTX6 U768 ( .A(n599), .B(n598), .Z(n1595) );
  ND2SVTX2 U769 ( .A(n1497), .B(n1498), .Z(n1493) );
  NR2SVTX2 U770 ( .A(n1535), .B(n445), .Z(n1540) );
  AO7SVTX2 U771 ( .A(n648), .B(n1500), .C(n1499), .Z(n649) );
  B_ND2SVTX2 U772 ( .A(n1582), .B(n334), .Z(n1583) );
  IVSVTX4 U773 ( .A(n447), .Z(n1502) );
  F_ND2SVTX1 U774 ( .A(n1734), .B(n1718), .Z(n1723) );
  OR2SVTX2 U775 ( .A(n1726), .B(n220), .Z(n1550) );
  ND2ASVTX4 U776 ( .A(n1446), .B(n670), .Z(n1745) );
  BFSVTX4 U777 ( .A(n1744), .Z(n443) );
  NR2SVTX4 U778 ( .A(n1417), .B(n1416), .Z(n1749) );
  AO2ABSVTX6 U779 ( .C(n873), .D(n767), .A(n875), .B(n252), .Z(n857) );
  IVSVTX2 U780 ( .A(n331), .Z(n688) );
  ND2SVTX4 U781 ( .A(n570), .B(n564), .Z(n563) );
  AO2SVTX4 U782 ( .A(n873), .B(n403), .C(n637), .D(n1420), .Z(n636) );
  NR3ABSVTX6 U783 ( .A(n253), .B(n654), .C(n1285), .Z(n689) );
  NR2SVTX4 U784 ( .A(n490), .B(n489), .Z(n1377) );
  ND2ASVTX4 U785 ( .A(n1238), .B(n1237), .Z(n1515) );
  ND2SVTX2 U786 ( .A(n223), .B(n1335), .Z(n489) );
  IVSVTX6 U787 ( .A(n1468), .Z(n237) );
  F_ND2ASVTX2 U788 ( .A(O[27]), .B(n1332), .Z(n1335) );
  MUX21NSVTX6 U789 ( .A(n826), .B(n276), .S(n766), .Z(n659) );
  IVSVTX6 U790 ( .A(n1252), .Z(n1275) );
  MUX21NSVTX4 U791 ( .A(n1392), .B(n1391), .S(n424), .Z(n1393) );
  ND2SVTX6 U792 ( .A(n285), .B(n231), .Z(n634) );
  ND2SVTX4 U793 ( .A(n1078), .B(n1079), .Z(n510) );
  MUX21NSVTX6 U794 ( .A(n1132), .B(n1158), .S(n871), .Z(n1396) );
  IVSVTX4 U795 ( .A(n1276), .Z(n765) );
  AO2SVTX4 U796 ( .A(n863), .B(n1219), .C(n862), .D(n1222), .Z(n861) );
  IVSVTX10 U797 ( .A(n593), .Z(n1184) );
  IVSVTX8 U798 ( .A(n540), .Z(n233) );
  IVSVTX8 U799 ( .A(n1224), .Z(n1203) );
  IVSVTX4 U800 ( .A(n719), .Z(n234) );
  AO2SVTX4 U801 ( .A(n243), .B(N[3]), .C(n469), .D(n666), .Z(n665) );
  CTIVSVTX2 U802 ( .A(n1060), .Z(n918) );
  IVSVTX4 U803 ( .A(N[3]), .Z(n1135) );
  IVSVTX6 U804 ( .A(N[21]), .Z(n1054) );
  AO7SVTX6 U805 ( .A(n630), .B(n626), .C(n624), .Z(n1615) );
  NR2SVTX6 U806 ( .A(n628), .B(n1568), .Z(n1643) );
  ND2SVTX6 U807 ( .A(n1523), .B(n452), .Z(n621) );
  ND2SVTX2 U808 ( .A(n465), .B(n1541), .Z(n464) );
  NR2SVTX2 U809 ( .A(n900), .B(n1542), .Z(n466) );
  AO7ASVTX4 U810 ( .A(n526), .B(n899), .C(n529), .Z(n531) );
  AO6SVTX2 U811 ( .A(n1550), .B(n526), .C(n530), .Z(n529) );
  B_ND2SVTX1 U812 ( .A(n327), .B(n436), .Z(n1656) );
  CTIVSVTX2 U813 ( .A(n327), .Z(n1690) );
  B_ND2SVTX2 U814 ( .A(n247), .B(n1657), .Z(n1659) );
  IVSVTX4 U815 ( .A(n1749), .Z(n1758) );
  B_ND2SVTX1 U816 ( .A(n686), .B(n1756), .Z(n1761) );
  AO7SVTX1 U817 ( .A(n1751), .B(n790), .C(n686), .Z(n1752) );
  IVSVTX2 U818 ( .A(n843), .Z(n842) );
  ND2ASVTX4 U819 ( .A(n1404), .B(n1447), .Z(n1744) );
  ND2SVTX4 U820 ( .A(n577), .B(n576), .Z(n843) );
  IVSVTX2 U821 ( .A(n525), .Z(n524) );
  B_ND2SVTX2 U822 ( .A(n1353), .B(n1547), .Z(n1520) );
  IVSVTX2 U823 ( .A(n844), .Z(n576) );
  ND2ASVTX6 U824 ( .A(n1248), .B(n1351), .Z(n523) );
  IVSVTX2 U825 ( .A(n1331), .Z(n413) );
  IVSVTX2 U826 ( .A(n1481), .Z(n559) );
  CTIVSVTX4 U827 ( .A(n1300), .Z(n1305) );
  IVSVTX4 U828 ( .A(n1475), .Z(n1331) );
  IVSVTX4 U829 ( .A(n875), .Z(n849) );
  BFSVTX4 U830 ( .A(n1299), .Z(n648) );
  NR2ASVTX4 U831 ( .A(n1451), .B(n875), .Z(n1438) );
  IVSVTX4 U832 ( .A(n1480), .Z(n567) );
  ND2SVTX6 U833 ( .A(n1082), .B(n1081), .Z(n1299) );
  IVSVTX2 U834 ( .A(n1377), .Z(n642) );
  IVSVTX6 U835 ( .A(n460), .Z(n236) );
  IVSVTX2 U836 ( .A(n1339), .Z(n1348) );
  IVSVTX10 U837 ( .A(n1184), .Z(n239) );
  ND3SVTX4 U838 ( .A(n815), .B(n1314), .C(n233), .Z(n1317) );
  IVSVTX12 U839 ( .A(n1186), .Z(n240) );
  IVSVTX2 U840 ( .A(n234), .Z(n717) );
  IVSVTX4 U841 ( .A(n428), .Z(n241) );
  IVSVTX4 U842 ( .A(n1222), .Z(n242) );
  ND2ASVTX6 U843 ( .A(n1218), .B(n1217), .Z(n1314) );
  IVSVTX2 U844 ( .A(n719), .Z(n747) );
  BFSVTX2 U845 ( .A(n959), .Z(O[31]) );
  ND4ABSVTX6 U846 ( .A(n955), .B(n956), .C(n954), .D(n260), .Z(n520) );
  IVSVTX4 U847 ( .A(n793), .Z(n796) );
  BFSVTX4 U848 ( .A(n479), .Z(n1136) );
  IVSVTX6 U849 ( .A(n1099), .Z(n398) );
  IVSVTX2 U850 ( .A(N[0]), .Z(n1137) );
  BFSVTX8 U851 ( .A(N[23]), .Z(n1099) );
  BFSVTX12 U852 ( .A(N[11]), .Z(n245) );
  B_ND2SVTX2 U853 ( .A(n1649), .B(n1648), .Z(n1650) );
  IVSVTX2 U854 ( .A(n630), .Z(n1621) );
  IVSVTX4 U855 ( .A(n1612), .Z(n1613) );
  F_AN2SVTX2 U856 ( .A(n1604), .B(n1603), .Z(n936) );
  NR2ASVTX8 U857 ( .A(n450), .B(n1587), .Z(n1638) );
  B_ND2SVTX2 U858 ( .A(n1625), .B(n931), .Z(n1626) );
  B_ND2SVTX2 U859 ( .A(n1494), .B(n1493), .Z(n1495) );
  AO7SVTX4 U860 ( .A(n1526), .B(n621), .C(n1525), .Z(n598) );
  ND2SVTX6 U861 ( .A(n1505), .B(n1504), .Z(n737) );
  NR2SVTX6 U862 ( .A(n477), .B(n940), .Z(n1651) );
  OR2SVTX2 U863 ( .A(n1624), .B(n1623), .Z(n931) );
  F_AN2SVTX2 U864 ( .A(n684), .B(n1513), .Z(n1566) );
  IVSVTX2 U865 ( .A(n466), .Z(n465) );
  B_ND2SVTX2 U866 ( .A(n526), .B(n527), .Z(n1662) );
  ND2SVTX6 U867 ( .A(n1553), .B(n531), .Z(n1565) );
  B_ND2SVTX2 U868 ( .A(n528), .B(n899), .Z(n527) );
  IVSVTX2 U869 ( .A(n625), .Z(n573) );
  AO6SVTX2 U870 ( .A(n1732), .B(n880), .C(n864), .Z(n1655) );
  B_ND2SVTX2 U871 ( .A(n1557), .B(n1559), .Z(n1562) );
  IVSVTX2 U872 ( .A(n1584), .Z(n625) );
  CTIVSVTX2 U873 ( .A(n449), .Z(n1538) );
  B_ND2SVTX2 U874 ( .A(n1661), .B(n1553), .Z(n1663) );
  NR2SVTX2 U875 ( .A(n902), .B(n1687), .Z(n1669) );
  B_ND2SVTX2 U876 ( .A(n1530), .B(n447), .Z(n1543) );
  AO7SVTX1 U877 ( .A(n1690), .B(n1689), .C(n436), .Z(n1691) );
  B_ND2SVTX2 U878 ( .A(n1556), .B(n1537), .Z(n1564) );
  B_ND2SVTX2 U879 ( .A(n1674), .B(n1677), .Z(n1680) );
  CTIVSVTX2 U880 ( .A(n1661), .Z(n530) );
  IVSVTX2 U881 ( .A(n1551), .Z(n526) );
  F_EOSVTX2 U882 ( .A(n1761), .B(n1760), .Z(O[0]) );
  AO7SVTX1 U883 ( .A(n462), .B(n1704), .C(n483), .Z(n1705) );
  IVSVTX6 U884 ( .A(n1479), .Z(n1675) );
  IVSVTX6 U885 ( .A(n439), .Z(n1291) );
  B_ND2SVTX2 U886 ( .A(n1710), .B(n483), .Z(n1715) );
  AO2ABSVTX4 U887 ( .C(n921), .D(n727), .A(n875), .B(n1301), .Z(n613) );
  IVSVTX4 U888 ( .A(n1242), .Z(n501) );
  NR2ASVTX6 U889 ( .A(n306), .B(n1307), .Z(n1726) );
  IVSVTX4 U890 ( .A(n1735), .Z(n1720) );
  ND2ASVTX6 U891 ( .A(n237), .B(n1472), .Z(n1701) );
  IVSVTX6 U892 ( .A(n1465), .Z(n1703) );
  ND2SVTX6 U893 ( .A(n643), .B(n1375), .Z(n574) );
  ND3ABSVTX4 U894 ( .A(n1300), .B(n335), .C(n1303), .Z(n727) );
  ND3ABSVTX6 U895 ( .A(n603), .B(n1443), .C(n444), .Z(n504) );
  NR2SVTX2 U896 ( .A(n790), .B(n1749), .Z(n1753) );
  ND2ASVTX4 U897 ( .A(n1406), .B(n842), .Z(n1415) );
  B_ND2SVTX1 U898 ( .A(n1748), .B(n1747), .Z(n1755) );
  NR2SVTX4 U899 ( .A(n1234), .B(n600), .Z(n503) );
  IVSVTX4 U900 ( .A(n585), .Z(n586) );
  ND3ASVTX6 U901 ( .A(n1248), .B(n286), .C(n699), .Z(n585) );
  ND2SVTX6 U902 ( .A(n802), .B(n696), .Z(n698) );
  ND2ASVTX4 U903 ( .A(n1468), .B(n1469), .Z(n525) );
  NR2SVTX4 U904 ( .A(n1301), .B(n1305), .Z(n676) );
  IVSVTX2 U905 ( .A(n1321), .Z(n646) );
  IVSVTX2 U906 ( .A(n1301), .Z(n335) );
  IVSVTX4 U907 ( .A(n710), .Z(n709) );
  IVSVTX4 U908 ( .A(n521), .Z(n248) );
  NR2ASVTX6 U909 ( .A(n1379), .B(n886), .Z(n584) );
  IVSVTX4 U910 ( .A(n875), .Z(n637) );
  IVSVTX6 U911 ( .A(n1379), .Z(n250) );
  IVSVTX2 U912 ( .A(n1510), .Z(n922) );
  NR2SVTX4 U913 ( .A(n491), .B(n1349), .Z(n488) );
  IVSVTX4 U914 ( .A(n616), .Z(n283) );
  IVSVTX4 U915 ( .A(n1446), .Z(n1404) );
  ND2SVTX4 U916 ( .A(n305), .B(n1193), .Z(n304) );
  CTIVSVTX6 U917 ( .A(n1574), .Z(n253) );
  NR3ABSVTX6 U918 ( .A(n1407), .B(n1310), .C(n735), .Z(n1354) );
  IVSVTX2 U919 ( .A(n1429), .Z(n653) );
  ND2SVTX4 U920 ( .A(n1214), .B(n1104), .Z(n1074) );
  ND2ASVTX4 U921 ( .A(n1183), .B(n1104), .Z(n1105) );
  IVSVTX2 U922 ( .A(n1400), .Z(n255) );
  ND3SVTX4 U923 ( .A(n1078), .B(n1079), .C(n231), .Z(n669) );
  IVSVTX2 U924 ( .A(n1272), .Z(n723) );
  IVSVTX8 U925 ( .A(n456), .Z(n887) );
  IVSVTX4 U926 ( .A(n806), .Z(n610) );
  AO7SVTX6 U927 ( .A(n1226), .B(n1225), .C(n596), .Z(n1262) );
  IVSVTX2 U928 ( .A(n317), .Z(n1385) );
  ND2SVTX6 U929 ( .A(n732), .B(n733), .Z(n730) );
  IVSVTX12 U930 ( .A(n266), .Z(n371) );
  AO6CSVTX6 U931 ( .A(n1056), .B(n1057), .C(n1280), .Z(n372) );
  IVSVTX2 U932 ( .A(n1413), .Z(n550) );
  IVSVTX4 U933 ( .A(n878), .Z(n1342) );
  ND2SVTX4 U934 ( .A(n352), .B(n351), .Z(n799) );
  IVSVTX2 U935 ( .A(n819), .Z(n823) );
  IVSVTX4 U936 ( .A(n1072), .Z(n850) );
  IVSVTX2 U937 ( .A(n1035), .Z(n303) );
  IVSVTX4 U938 ( .A(n718), .Z(n715) );
  IVSVTX2 U939 ( .A(n882), .Z(n788) );
  NR2SVTX2 U940 ( .A(n1007), .B(n1006), .Z(n752) );
  IVSVTX2 U941 ( .A(n1187), .Z(n879) );
  NR2SVTX4 U942 ( .A(n1280), .B(n1215), .Z(n725) );
  IVSVTX4 U943 ( .A(n896), .Z(n1200) );
  ND3SVTX8 U944 ( .A(n1022), .B(n406), .C(n405), .Z(n354) );
  IVSVTX4 U945 ( .A(n1388), .Z(n257) );
  IVSVTX2 U946 ( .A(n1031), .Z(n1033) );
  IVSVTX2 U947 ( .A(n308), .Z(n307) );
  IVSVTX2 U948 ( .A(n1139), .Z(n333) );
  IVSVTX12 U949 ( .A(n519), .Z(n258) );
  CTIVSVTX4 U950 ( .A(n292), .Z(n291) );
  AO7SVTX6 U951 ( .A(n944), .B(n796), .C(n1010), .Z(n821) );
  ND2SVTX4 U952 ( .A(n987), .B(n986), .Z(n1150) );
  IVSVTX8 U953 ( .A(n1009), .Z(n594) );
  IVSVTX8 U954 ( .A(n473), .Z(n912) );
  IVSVTX2 U955 ( .A(n1025), .Z(n430) );
  IVSVTX4 U956 ( .A(n394), .Z(n393) );
  IVSVTX4 U957 ( .A(n975), .Z(n606) );
  CTIVSVTX2 U958 ( .A(n1001), .Z(n1002) );
  IVSVTX8 U959 ( .A(n363), .Z(n260) );
  ND2SVTX6 U960 ( .A(n475), .B(n971), .Z(n380) );
  BFSVTX4 U961 ( .A(N[19]), .Z(n469) );
  IVSVTX8 U962 ( .A(N[26]), .Z(n1023) );
  NR2SVTX6 U963 ( .A(N[8]), .B(N[11]), .Z(n794) );
  IVSVTX6 U964 ( .A(N[12]), .Z(n263) );
  IVSVTX6 U965 ( .A(N[31]), .Z(n264) );
  ND4ABSVTX8 U966 ( .A(n251), .B(n1360), .C(n708), .D(n568), .Z(n720) );
  ND2SVTX4 U967 ( .A(n810), .B(n265), .Z(n1182) );
  IVSVTX4 U968 ( .A(n1262), .Z(n265) );
  IVSVTX4 U969 ( .A(n267), .Z(n320) );
  ND2SVTX4 U970 ( .A(n401), .B(n728), .Z(n267) );
  ND2ASVTX8 U971 ( .A(n1401), .B(n729), .Z(n728) );
  IVSVTX4 U972 ( .A(n270), .Z(n729) );
  ND2ASVTX8 U973 ( .A(n1113), .B(n924), .Z(n1401) );
  AO6ABSVTX6 U974 ( .A(n358), .B(n788), .C(n268), .Z(n401) );
  IVSVTX4 U975 ( .A(n402), .Z(n268) );
  ND2SVTX6 U976 ( .A(n887), .B(n759), .Z(n269) );
  IVSVTX4 U977 ( .A(n1401), .Z(n274) );
  ND2SVTX4 U978 ( .A(n753), .B(n271), .Z(n270) );
  ND3ASVTX6 U979 ( .A(n259), .B(n753), .C(n271), .Z(n273) );
  ND2SVTX6 U980 ( .A(n414), .B(n273), .Z(n456) );
  ND2ASVTX8 U981 ( .A(n275), .B(n659), .Z(n1574) );
  ND4ABSVTX8 U982 ( .A(n276), .B(n275), .C(n1110), .D(n433), .Z(n432) );
  ND2SVTX4 U983 ( .A(n424), .B(n276), .Z(n660) );
  ND3SVTX6 U984 ( .A(n780), .B(n779), .C(n781), .Z(n276) );
  CTIVSVTX6 U985 ( .A(n1452), .Z(n279) );
  AO6ASVTX8 U986 ( .A(n1744), .B(n1740), .C(n277), .Z(n1719) );
  IVSVTX4 U987 ( .A(n1739), .Z(n277) );
  ND2ASVTX8 U988 ( .A(n754), .B(n278), .Z(n1740) );
  IVSVTX4 U989 ( .A(n1448), .Z(n278) );
  ND2SVTX4 U990 ( .A(n1445), .B(n1444), .Z(n1447) );
  AO7SVTX8 U991 ( .A(n1455), .B(n1719), .C(n280), .Z(n1456) );
  AO6SVTX8 U992 ( .A(n1720), .B(n1716), .C(n281), .Z(n280) );
  ND2SVTX6 U993 ( .A(n1734), .B(n1716), .Z(n1455) );
  ND2ASVTX6 U994 ( .A(n255), .B(n282), .Z(n1734) );
  IVSVTX4 U995 ( .A(n1450), .Z(n282) );
  AN2SVTX8 U996 ( .A(n284), .B(n283), .Z(n615) );
  ND2SVTX4 U997 ( .A(n766), .B(n285), .Z(n284) );
  AO7SVTX8 U998 ( .A(n1285), .B(n801), .C(n1519), .Z(n286) );
  IVSVTX4 U999 ( .A(n287), .Z(n1657) );
  AO20SVTX8 U1000 ( .A(n1353), .B(n318), .C(n857), .D(n250), .Z(n287) );
  IVSVTX10 U1001 ( .A(n288), .Z(n830) );
  ND3ABSVTX6 U1002 ( .A(n814), .B(n1041), .C(n870), .Z(n288) );
  ND2SVTX4 U1003 ( .A(n1219), .B(n830), .Z(n1254) );
  ND2ASVTX8 U1004 ( .A(n288), .B(n1213), .Z(n712) );
  ND2SVTX4 U1005 ( .A(n830), .B(n785), .Z(n837) );
  NR2SVTX6 U1006 ( .A(N[31]), .B(N[28]), .Z(n370) );
  ND3SVTX4 U1007 ( .A(n605), .B(n289), .C(n1249), .Z(n846) );
  IVSVTX4 U1008 ( .A(n290), .Z(n745) );
  ND2SVTX4 U1009 ( .A(n1390), .B(n290), .Z(n1256) );
  MUX21NSVTX6 U1010 ( .A(n1252), .B(n290), .S(n428), .Z(n1364) );
  ND3SVTX8 U1011 ( .A(n713), .B(n712), .C(n711), .Z(n290) );
  ND2ASVTX8 U1012 ( .A(n357), .B(n1113), .Z(n293) );
  AO7ABSVTX4 U1013 ( .A(n293), .B(n409), .C(n749), .Z(n1127) );
  AO8ASVTX6 U1014 ( .A(n361), .B(n1116), .C(n1175), .D(n1157), .Z(n1121) );
  NR2ASVTX8 U1015 ( .A(n291), .B(n293), .Z(n1157) );
  NR2SVTX8 U1016 ( .A(n1115), .B(n1172), .Z(n292) );
  ND2SVTX8 U1017 ( .A(n507), .B(n508), .Z(n1245) );
  ND4SVTX4 U1018 ( .A(n507), .B(n1082), .C(n508), .D(n1081), .Z(n1300) );
  AO2SVTX8 U1019 ( .A(n731), .B(n1129), .C(n1134), .D(N[3]), .Z(n294) );
  NR2ASVTX8 U1020 ( .A(n734), .B(n294), .Z(n1384) );
  ND2SVTX8 U1021 ( .A(n1426), .B(n1424), .Z(n1433) );
  NR2SVTX6 U1022 ( .A(n295), .B(n296), .Z(n400) );
  ND2ASVTX8 U1023 ( .A(n296), .B(n898), .Z(n1420) );
  IVSVTX6 U1024 ( .A(n1257), .Z(n1282) );
  AO6SVTX8 U1025 ( .A(n329), .B(n480), .C(n1259), .Z(n1365) );
  MUX21NSVTX8 U1026 ( .A(n1121), .B(n1126), .S(n421), .Z(n1397) );
  IVSVTX8 U1027 ( .A(n869), .Z(n870) );
  ND2SVTX4 U1028 ( .A(n240), .B(n1077), .Z(n1065) );
  ND2SVTX4 U1029 ( .A(n766), .B(n1080), .Z(n668) );
  IVSVTX4 U1030 ( .A(n1051), .Z(n297) );
  ND3SVTX6 U1031 ( .A(n1085), .B(n1172), .C(n1084), .Z(n298) );
  IVSVTX10 U1032 ( .A(n1134), .Z(n731) );
  ENSVTX8 U1033 ( .A(n1475), .B(n299), .Z(n639) );
  ND4SVTX6 U1034 ( .A(n237), .B(n348), .C(n236), .D(n1398), .Z(n299) );
  ND2SVTX4 U1035 ( .A(n379), .B(n407), .Z(n406) );
  IVSVTX4 U1036 ( .A(n358), .Z(n1251) );
  IVSVTX4 U1037 ( .A(n870), .Z(n332) );
  IVSVTX4 U1038 ( .A(n682), .Z(n663) );
  ND3ABSVTX8 U1039 ( .A(n893), .B(n947), .C(n301), .Z(n1143) );
  IVSVTX4 U1040 ( .A(n895), .Z(n301) );
  AO17ASVTX8 U1041 ( .A(n1406), .B(n874), .C(n549), .D(n1412), .Z(n548) );
  ND3ABSVTX8 U1042 ( .A(n303), .B(n1050), .C(n935), .Z(n387) );
  NR2SVTX4 U1043 ( .A(n304), .B(n1260), .Z(n760) );
  NR2SVTX4 U1044 ( .A(n1258), .B(n1194), .Z(n305) );
  IVSVTX10 U1045 ( .A(n385), .Z(n924) );
  AO4ABSVTX6 U1046 ( .C(n1443), .D(n1417), .A(n1406), .B(n249), .Z(n549) );
  NR2SVTX4 U1047 ( .A(n306), .B(n1480), .Z(n557) );
  NR2SVTX4 U1048 ( .A(n823), .B(n1180), .Z(n319) );
  IVSVTX6 U1049 ( .A(n1140), .Z(n759) );
  AO3ASVTX6 U1050 ( .A(n371), .B(n838), .C(n968), .D(n969), .Z(n533) );
  ND2SVTX4 U1051 ( .A(n1180), .B(n1179), .Z(n359) );
  AO7SVTX6 U1052 ( .A(n361), .B(n1155), .C(n307), .Z(n1179) );
  NR2SVTX4 U1053 ( .A(n360), .B(n1154), .Z(n308) );
  IVSVTX4 U1054 ( .A(n1343), .Z(n309) );
  BFSVTX2 U1055 ( .A(n1736), .Z(n310) );
  IVSVTX4 U1056 ( .A(n1317), .Z(n1340) );
  NR2ASVTX6 U1057 ( .A(n1449), .B(n875), .Z(n1440) );
  IVSVTX6 U1058 ( .A(n748), .Z(n421) );
  ND3ASVTX8 U1059 ( .A(n1428), .B(n458), .C(n1430), .Z(n1450) );
  NR2SVTX4 U1060 ( .A(n218), .B(n682), .Z(n1006) );
  ND2SVTX6 U1061 ( .A(n342), .B(n912), .Z(n349) );
  IVSVTX4 U1062 ( .A(n349), .Z(n357) );
  IVSVTX8 U1063 ( .A(n1154), .Z(n1113) );
  IVSVTX12 U1064 ( .A(n814), .Z(n815) );
  AO4SVTX8 U1065 ( .A(n1215), .B(n382), .C(n1223), .D(n641), .Z(n336) );
  ND4SVTX6 U1066 ( .A(n1350), .B(n312), .C(n311), .D(n488), .Z(n487) );
  IVSVTX4 U1067 ( .A(n492), .Z(n311) );
  IVSVTX4 U1068 ( .A(n313), .Z(n312) );
  ND2SVTX4 U1069 ( .A(n314), .B(n1347), .Z(n313) );
  IVSVTX4 U1070 ( .A(n1141), .Z(n314) );
  ND2SVTX4 U1071 ( .A(n315), .B(n806), .Z(n1339) );
  ND3SVTX6 U1072 ( .A(n1325), .B(n435), .C(n428), .Z(n315) );
  ND2SVTX4 U1073 ( .A(n1324), .B(n485), .Z(n1343) );
  ND2ASVTX8 U1074 ( .A(n241), .B(n1329), .Z(n339) );
  AO6SVTX6 U1075 ( .A(n1403), .B(n378), .C(n377), .Z(n376) );
  AO7SVTX8 U1076 ( .A(n1248), .B(n1405), .C(n376), .Z(n1418) );
  ND3SVTX8 U1077 ( .A(n1150), .B(n235), .C(n353), .Z(n998) );
  IVSVTX4 U1078 ( .A(n1709), .Z(n522) );
  ND2ASVTX8 U1079 ( .A(n316), .B(n338), .Z(n1709) );
  ENSVTX8 U1080 ( .A(n322), .B(n858), .Z(n318) );
  ND2SVTX6 U1081 ( .A(n1094), .B(n240), .Z(n1091) );
  ND2ASVTX8 U1082 ( .A(n1248), .B(n1359), .Z(n726) );
  ND2SVTX6 U1083 ( .A(n238), .B(n852), .Z(n1702) );
  NR3ABSVTX2 U1084 ( .A(n754), .B(n1230), .C(n1047), .Z(n644) );
  NR2SVTX4 U1085 ( .A(n263), .B(n999), .Z(n1061) );
  AO2SVTX4 U1086 ( .A(n1431), .B(n874), .C(n249), .D(n1461), .Z(n1432) );
  ND2ASVTX8 U1087 ( .A(n1453), .B(n1452), .Z(n1454) );
  NR2ASVTX6 U1088 ( .A(n386), .B(n1152), .Z(n853) );
  ND3SVTX6 U1089 ( .A(n606), .B(n260), .C(n607), .Z(n386) );
  AO7ABSVTX8 U1090 ( .A(N[5]), .B(n1038), .C(n777), .Z(n914) );
  ND3SVTX8 U1091 ( .A(n371), .B(n1390), .C(n903), .Z(n806) );
  ND3SVTX6 U1092 ( .A(n358), .B(n1170), .C(n319), .Z(n498) );
  ND2SVTX4 U1093 ( .A(n1224), .B(n1208), .Z(n1324) );
  ND4SVTX4 U1094 ( .A(n400), .B(n366), .C(n399), .D(n320), .Z(n735) );
  ND2SVTX4 U1095 ( .A(n1189), .B(n321), .Z(n1217) );
  IVSVTX4 U1096 ( .A(n258), .Z(n321) );
  BFSVTX1 U1097 ( .A(n1293), .Z(n322) );
  ND3ABSVTX8 U1098 ( .A(n1284), .B(n1283), .C(n1282), .Z(n1379) );
  ND3SVTX8 U1099 ( .A(n344), .B(n1254), .C(n1253), .Z(n1268) );
  IVSVTX8 U1100 ( .A(N[28]), .Z(n828) );
  IVSVTX8 U1101 ( .A(n323), .Z(n1273) );
  AO7SVTX8 U1102 ( .A(n231), .B(n1220), .C(n745), .Z(n744) );
  IVSVTX6 U1103 ( .A(n924), .Z(n1224) );
  ND3SVTX8 U1104 ( .A(n606), .B(n607), .C(n260), .Z(n608) );
  ND2SVTX4 U1105 ( .A(n1192), .B(n835), .Z(n323) );
  NR3SVTX8 U1106 ( .A(n638), .B(n325), .C(n324), .Z(n1264) );
  NR2SVTX4 U1107 ( .A(n1181), .B(n1262), .Z(n324) );
  ND2SVTX4 U1108 ( .A(n1263), .B(n498), .Z(n325) );
  IVSVTX10 U1109 ( .A(n371), .Z(n1221) );
  NR3SVTX8 U1110 ( .A(n1259), .B(n746), .C(n744), .Z(n1227) );
  IVSVTX6 U1111 ( .A(N[29]), .Z(n453) );
  ND2ASVTX8 U1112 ( .A(N[4]), .B(n1053), .Z(n990) );
  IVSVTX8 U1113 ( .A(n1369), .Z(n568) );
  ND2SVTX8 U1114 ( .A(n930), .B(n1587), .Z(n1639) );
  NR2SVTX8 U1115 ( .A(n976), .B(n446), .Z(n607) );
  ENSVTX6 U1116 ( .A(n1427), .B(n854), .Z(n1431) );
  IVSVTX8 U1117 ( .A(n1213), .Z(n1107) );
  IVSVTX10 U1118 ( .A(n371), .Z(n871) );
  ND3SVTX8 U1119 ( .A(n395), .B(n390), .C(n330), .Z(n355) );
  AO17SVTX8 U1120 ( .A(n393), .B(n388), .C(n389), .D(n260), .Z(n330) );
  ND3ABSVTX8 U1121 ( .A(n333), .B(n332), .C(n415), .Z(n414) );
  IVSVTX6 U1122 ( .A(n786), .Z(n1004) );
  ND3SVTX8 U1123 ( .A(n472), .B(n471), .C(n441), .Z(n364) );
  AO7SVTX8 U1124 ( .A(n1045), .B(n1080), .C(n615), .Z(n1498) );
  IVSVTX12 U1125 ( .A(n641), .Z(n891) );
  IVSVTX12 U1126 ( .A(n595), .Z(n999) );
  ND3SVTX8 U1127 ( .A(n1364), .B(n1282), .C(n1368), .Z(n710) );
  ND2ASVTX8 U1128 ( .A(n1030), .B(n437), .Z(n1024) );
  IVSVTX8 U1129 ( .A(n1114), .Z(n1084) );
  BFSVTX1 U1130 ( .A(n353), .Z(n337) );
  AO7SVTX8 U1131 ( .A(n1353), .B(n639), .C(n467), .Z(n338) );
  IVSVTX4 U1132 ( .A(n338), .Z(n852) );
  AO3ASVTX6 U1133 ( .A(n424), .B(n1323), .C(n339), .D(n1342), .Z(n460) );
  ND2ASVTX8 U1134 ( .A(n340), .B(n309), .Z(n1329) );
  IVSVTX4 U1135 ( .A(n1341), .Z(n340) );
  ND2SVTX8 U1136 ( .A(n1054), .B(n1058), .Z(n422) );
  IVSVTX6 U1137 ( .A(N[20]), .Z(n1058) );
  NR2SVTX4 U1138 ( .A(n1027), .B(n342), .Z(n407) );
  ND3ASVTX6 U1139 ( .A(N[22]), .B(n398), .C(n244), .Z(n342) );
  NR2SVTX6 U1140 ( .A(n343), .B(n514), .Z(n1193) );
  ND3SVTX8 U1141 ( .A(n326), .B(n516), .C(n344), .Z(n343) );
  ND2SVTX8 U1142 ( .A(n891), .B(n345), .Z(n344) );
  ND2SVTX6 U1143 ( .A(n346), .B(n347), .Z(n473) );
  NR2SVTX6 U1144 ( .A(N[24]), .B(N[26]), .Z(n347) );
  ND3SVTX8 U1145 ( .A(n348), .B(n237), .C(n1398), .Z(n429) );
  ND2SVTX4 U1146 ( .A(n946), .B(n349), .Z(n820) );
  NR2SVTX4 U1147 ( .A(n1174), .B(n385), .Z(n351) );
  AO17ASVTX4 U1148 ( .A(n1173), .B(n1172), .C(n1171), .D(n815), .Z(n352) );
  ND2SVTX8 U1149 ( .A(n988), .B(n379), .Z(n353) );
  IVSVTX4 U1150 ( .A(n354), .Z(n1187) );
  ND2ASVTX8 U1151 ( .A(n354), .B(n1133), .Z(n1134) );
  NR2SVTX4 U1152 ( .A(n354), .B(n355), .Z(n408) );
  IVSVTX10 U1153 ( .A(n355), .Z(n1133) );
  ND2SVTX8 U1154 ( .A(n356), .B(n1354), .Z(n1369) );
  ND4SVTX4 U1155 ( .A(n1363), .B(n356), .C(n1365), .D(n1354), .Z(n571) );
  IVSVTX12 U1156 ( .A(n423), .Z(n358) );
  ND2SVTX4 U1157 ( .A(n358), .B(n359), .Z(n596) );
  IVSVTX4 U1158 ( .A(n423), .Z(n892) );
  ND3ABSVTX8 U1159 ( .A(n1265), .B(n1437), .C(n1264), .Z(n362) );
  ND3SVTX8 U1160 ( .A(n953), .B(n609), .C(n952), .Z(n363) );
  NR3SVTX8 U1161 ( .A(n1014), .B(n363), .C(n446), .Z(n391) );
  ND2SVTX4 U1162 ( .A(n424), .B(n364), .Z(n1095) );
  ND2SVTX4 U1163 ( .A(O[27]), .B(n364), .Z(n656) );
  ND2ASVTX8 U1164 ( .A(n1143), .B(n520), .Z(n365) );
  IVSVTX10 U1165 ( .A(n365), .Z(n519) );
  ND2SVTX4 U1166 ( .A(n776), .B(n365), .Z(n1069) );
  ND3SVTX8 U1167 ( .A(n401), .B(n366), .C(n400), .Z(n1312) );
  ND2SVTX4 U1168 ( .A(n366), .B(n1393), .Z(n1446) );
  ND2SVTX8 U1169 ( .A(n1221), .B(n1131), .Z(n366) );
  ND2SVTX4 U1170 ( .A(n957), .B(n368), .Z(n976) );
  ND4ASVTX6 U1171 ( .A(N[27]), .B(n369), .C(n368), .D(n475), .Z(n394) );
  IVSVTX4 U1172 ( .A(N[16]), .Z(n958) );
  ND2SVTX8 U1173 ( .A(n370), .B(n1023), .Z(n446) );
  NR3ABSVTX8 U1174 ( .A(n661), .B(n662), .C(n372), .Z(n838) );
  NR2ASVTX8 U1175 ( .A(n403), .B(n375), .Z(n404) );
  ND3ASVTX8 U1176 ( .A(n644), .B(n374), .C(n373), .Z(n375) );
  ND2SVTX8 U1177 ( .A(n1577), .B(n1441), .Z(n373) );
  AO7SVTX6 U1178 ( .A(n687), .B(n404), .C(n1747), .Z(n476) );
  ND2SVTX4 U1179 ( .A(n1420), .B(n375), .Z(n1747) );
  ND2ASVTX8 U1180 ( .A(n256), .B(n1418), .Z(n687) );
  F_ENSVTX2 U1181 ( .A(n1446), .B(n1395), .Z(n1405) );
  ND2ASVTX8 U1182 ( .A(n638), .B(n582), .Z(n1461) );
  AO6SVTX4 U1183 ( .A(n397), .B(n379), .C(n396), .Z(n395) );
  NR2SVTX8 U1184 ( .A(n380), .B(n972), .Z(n379) );
  NR2SVTX4 U1185 ( .A(n815), .B(n385), .Z(n383) );
  ND2ASVTX8 U1186 ( .A(n815), .B(n266), .Z(n641) );
  ND2SVTX8 U1187 ( .A(n1205), .B(n1133), .Z(n385) );
  IVSVTX4 U1188 ( .A(n386), .Z(n776) );
  NR2SVTX4 U1189 ( .A(n1195), .B(n853), .Z(n1155) );
  NR2ASVTX6 U1190 ( .A(n1151), .B(n1172), .Z(n1195) );
  ND3SVTX8 U1191 ( .A(n371), .B(n1037), .C(n387), .Z(n1044) );
  NR3SVTX8 U1192 ( .A(n992), .B(n446), .C(n974), .Z(n388) );
  AO7SVTX8 U1193 ( .A(n957), .B(n972), .C(n264), .Z(n396) );
  CTIVSVTX4 U1194 ( .A(n1312), .Z(n434) );
  NR3SVTX8 U1195 ( .A(n730), .B(n1384), .C(n1386), .Z(n399) );
  NR2SVTX6 U1196 ( .A(n404), .B(n789), .Z(n1421) );
  ND2SVTX6 U1197 ( .A(n890), .B(n474), .Z(n405) );
  MUX21NSVTX8 U1198 ( .A(n1125), .B(n1127), .S(n748), .Z(n1130) );
  NR3ABSVTX8 U1199 ( .A(n759), .B(n887), .C(n1312), .Z(n1424) );
  ND2SVTX8 U1200 ( .A(n562), .B(n561), .Z(n410) );
  ND2SVTX8 U1201 ( .A(n559), .B(n410), .Z(n1672) );
  ND3SVTX4 U1202 ( .A(N[3]), .B(n1154), .C(n1205), .Z(n1389) );
  NR2SVTX6 U1203 ( .A(N[26]), .B(N[25]), .Z(n971) );
  IVSVTX4 U1204 ( .A(n411), .Z(n1471) );
  NR2SVTX4 U1205 ( .A(n884), .B(n639), .Z(n411) );
  ND2SVTX4 U1206 ( .A(n1311), .B(n1310), .Z(n418) );
  ND3SVTX8 U1207 ( .A(n1092), .B(n419), .C(n1091), .Z(n783) );
  AO7SVTX8 U1208 ( .A(n1478), .B(n1688), .C(n1685), .Z(n1479) );
  AO7SVTX8 U1209 ( .A(n454), .B(n455), .C(n413), .Z(n1685) );
  BFSVTX2 U1210 ( .A(N[13]), .Z(n1188) );
  IVSVTX6 U1211 ( .A(n519), .Z(n682) );
  ND2SVTX4 U1212 ( .A(n1084), .B(n416), .Z(n1197) );
  NR2SVTX4 U1213 ( .A(n1135), .B(n493), .Z(n416) );
  IVSVTX6 U1214 ( .A(n836), .Z(n874) );
  ND2ASVTX8 U1215 ( .A(n836), .B(n1376), .Z(n643) );
  IVSVTX12 U1216 ( .A(n358), .Z(n1411) );
  ND3SVTX6 U1217 ( .A(n1469), .B(n1470), .C(n1471), .Z(n1472) );
  BFSVTX6 U1218 ( .A(n1047), .Z(n417) );
  IVSVTX8 U1219 ( .A(n440), .Z(n595) );
  IVSVTX6 U1220 ( .A(n639), .Z(n1351) );
  AO5SVTX6 U1221 ( .A(n550), .B(n548), .C(n546), .Z(n1414) );
  ENSVTX6 U1222 ( .A(n1419), .B(n1407), .Z(n1410) );
  ND3ABSVTX8 U1223 ( .A(n1461), .B(n418), .C(n1398), .Z(n1313) );
  ND3ASVTX6 U1224 ( .A(n730), .B(n728), .C(n887), .Z(n757) );
  AO7ASVTX8 U1225 ( .A(n334), .B(n619), .C(n1582), .Z(n484) );
  IVSVTX4 U1226 ( .A(n425), .Z(n1363) );
  ND2ASVTX8 U1227 ( .A(n425), .B(n1365), .Z(n1360) );
  ND2ASVTX8 U1228 ( .A(n1373), .B(n554), .Z(n556) );
  ND2SVTX4 U1229 ( .A(n1745), .B(n1740), .Z(n1736) );
  ND3ASVTX6 U1230 ( .A(n815), .B(n1213), .C(n233), .Z(n419) );
  AO1SVTX4 U1231 ( .A(N[0]), .B(n1172), .C(n1176), .D(n361), .Z(n1156) );
  ND3SVTX8 U1232 ( .A(n1028), .B(n1187), .C(n1133), .Z(n423) );
  IVSVTX6 U1233 ( .A(n1378), .Z(n1664) );
  NR3ABSVTX2 U1234 ( .A(N[3]), .B(n1136), .C(n428), .Z(n867) );
  ENSVTX6 U1235 ( .A(n1631), .B(n1630), .Z(O[21]) );
  IVSVTX4 U1236 ( .A(n1133), .Z(n869) );
  AN2SVTX4 U1237 ( .A(n1379), .B(n1368), .Z(n928) );
  NR2SVTX8 U1238 ( .A(n807), .B(n1296), .Z(n1533) );
  BFSVTX4 U1239 ( .A(n1394), .Z(n426) );
  AO2SVTX6 U1240 ( .A(n731), .B(N[0]), .C(n1134), .D(N[1]), .Z(n1408) );
  AO2ABSVTX8 U1241 ( .C(n873), .D(n1355), .A(n1377), .B(n534), .Z(n1356) );
  NR2SVTX4 U1242 ( .A(n912), .B(n1117), .Z(n1145) );
  IVSVTX4 U1243 ( .A(n1114), .Z(n959) );
  IVSVTX2 U1244 ( .A(n1197), .Z(n1160) );
  ENSVTX8 U1245 ( .A(n236), .B(n429), .Z(n1352) );
  IVSVTX4 U1246 ( .A(n1258), .Z(n835) );
  AO7ASVTX8 U1247 ( .A(n430), .B(n1153), .C(n1024), .Z(n474) );
  NR3ABSVTX8 U1248 ( .A(n925), .B(n1111), .C(n432), .Z(n1112) );
  IVSVTX4 U1249 ( .A(n1238), .Z(n433) );
  ND3SVTX8 U1250 ( .A(n1208), .B(n859), .C(n1411), .Z(n1333) );
  ND2ASVTX8 U1251 ( .A(n1574), .B(n654), .Z(n697) );
  ND2SVTX8 U1252 ( .A(n558), .B(n556), .Z(n1376) );
  ND2SVTX6 U1253 ( .A(n928), .B(n1367), .Z(n832) );
  ND3SVTX8 U1254 ( .A(n1310), .B(n434), .C(n1394), .Z(n1229) );
  ND3SVTX8 U1255 ( .A(n694), .B(n693), .C(n692), .Z(n826) );
  ND2SVTX6 U1256 ( .A(n1700), .B(n522), .Z(n1473) );
  BFSVTX6 U1257 ( .A(N[9]), .Z(n438) );
  ND3SVTX6 U1258 ( .A(n798), .B(n252), .C(n797), .Z(n439) );
  ND2SVTX4 U1259 ( .A(n1084), .B(n519), .Z(n440) );
  ND2SVTX4 U1260 ( .A(n240), .B(n914), .Z(n441) );
  OR2SVTX8 U1261 ( .A(n856), .B(n1293), .Z(n1285) );
  AO7ABSVTX4 U1262 ( .A(n1093), .B(n486), .C(n617), .Z(n616) );
  BFSVTX4 U1263 ( .A(n1719), .Z(n442) );
  ENSVTX8 U1264 ( .A(n1453), .B(n755), .Z(n1442) );
  ND2ASVTX8 U1265 ( .A(n1443), .B(n1442), .Z(n1444) );
  AO5SVTX4 U1266 ( .A(n627), .B(n1651), .C(n1567), .Z(n1569) );
  AO6CSVTX8 U1267 ( .A(n741), .B(n675), .C(n1577), .Z(n679) );
  ND3SVTX8 U1268 ( .A(n1311), .B(n825), .C(n1182), .Z(n866) );
  IVSVTX4 U1269 ( .A(n602), .Z(n444) );
  ND2SVTX4 U1270 ( .A(n742), .B(n1228), .Z(n602) );
  BFSVTX1 U1271 ( .A(n1534), .Z(n445) );
  IVSVTX4 U1272 ( .A(n1578), .Z(n623) );
  ND3SVTX8 U1273 ( .A(n504), .B(n505), .C(n503), .Z(n1506) );
  ND2ASVTX8 U1274 ( .A(n805), .B(n709), .Z(n722) );
  IVSVTX8 U1275 ( .A(n608), .Z(n1114) );
  NR2SVTX4 U1276 ( .A(n747), .B(n266), .Z(n862) );
  ND3ASVTX8 U1277 ( .A(n676), .B(n679), .C(n680), .Z(n502) );
  ND3ASVTX8 U1278 ( .A(n1039), .B(n946), .C(n912), .Z(n800) );
  ND3SVTX4 U1279 ( .A(N[5]), .B(n1146), .C(n1016), .Z(n1011) );
  IVSVTX4 U1280 ( .A(n930), .Z(n450) );
  AO7SVTX4 U1281 ( .A(n1642), .B(n1638), .C(n901), .Z(n1636) );
  ND2SVTX6 U1282 ( .A(n984), .B(n983), .Z(n985) );
  IVSVTX4 U1283 ( .A(n496), .Z(n622) );
  ND3SVTX8 U1284 ( .A(n569), .B(n557), .C(n568), .Z(n558) );
  ND2SVTX4 U1285 ( .A(n563), .B(n565), .Z(n454) );
  ND3SVTX8 U1286 ( .A(n1439), .B(n833), .C(n834), .Z(n1448) );
  AO6SVTX8 U1287 ( .A(n1558), .B(n845), .C(n1298), .Z(n538) );
  BFSVTX1 U1288 ( .A(n1516), .Z(n457) );
  ENSVTX6 U1289 ( .A(n905), .B(n484), .Z(n1509) );
  ND2SVTX4 U1290 ( .A(n921), .B(n1431), .Z(n458) );
  MUX21NSVTX8 U1291 ( .A(n459), .B(n1179), .S(n748), .Z(n1164) );
  NR2SVTX4 U1292 ( .A(n1157), .B(n1156), .Z(n459) );
  IVSVTX2 U1293 ( .A(n1216), .Z(n1218) );
  ND2ASVTX8 U1294 ( .A(n1361), .B(n1364), .Z(n1373) );
  IVSVTX8 U1295 ( .A(n743), .Z(n740) );
  ND2ASVTX8 U1296 ( .A(n743), .B(n689), .Z(n589) );
  IVSVTX8 U1297 ( .A(n1250), .Z(n588) );
  IVSVTX10 U1298 ( .A(n1606), .Z(n1631) );
  NR2ASVTX8 U1299 ( .A(n371), .B(n1164), .Z(n638) );
  NR2SVTX8 U1300 ( .A(N[16]), .B(N[24]), .Z(n980) );
  ND3SVTX8 U1301 ( .A(n224), .B(n751), .C(n750), .Z(n1459) );
  AO17SVTX4 U1302 ( .A(n766), .B(n1267), .C(n1266), .D(n1276), .Z(n1272) );
  BFSVTX1 U1303 ( .A(n1573), .Z(n463) );
  F_ENSVTX2 U1304 ( .A(n1543), .B(n464), .Z(n1544) );
  AO2ABSVTX8 U1305 ( .C(n873), .D(n1352), .A(n236), .B(n534), .Z(n467) );
  ND2SVTX4 U1306 ( .A(n1219), .B(n891), .Z(n472) );
  ND2SVTX4 U1307 ( .A(n1546), .B(n1521), .Z(n1512) );
  AO7SVTX8 U1308 ( .A(n1601), .B(n1606), .C(n1600), .Z(n1627) );
  F_ND2ASVTX2 U1309 ( .A(n937), .B(n1627), .Z(n908) );
  EO3SVTX8 U1310 ( .A(n1572), .B(n771), .C(n629), .Z(n628) );
  IVSVTX8 U1311 ( .A(n695), .Z(n742) );
  ND2ASVTX8 U1312 ( .A(n695), .B(n740), .Z(n583) );
  ND3SVTX8 U1313 ( .A(n622), .B(n1509), .C(n1521), .Z(n604) );
  AO5NSVTX4 U1314 ( .A(n1584), .B(n572), .C(n581), .Z(n1589) );
  CTBUFSVTX8 U1315 ( .A(n633), .Z(n477) );
  AO7SVTX8 U1316 ( .A(n1728), .B(n220), .C(n1657), .Z(n1551) );
  IVSVTX8 U1317 ( .A(N[30]), .Z(n945) );
  AO8SVTX6 U1318 ( .A(n704), .B(n216), .C(n703), .D(n784), .Z(n702) );
  AO17CSVTX8 U1319 ( .A(n706), .B(n705), .C(n921), .D(n702), .Z(n839) );
  IVSVTX8 U1320 ( .A(n756), .Z(n1249) );
  BFSVTX1 U1321 ( .A(n893), .Z(n479) );
  AO7SVTX8 U1322 ( .A(n620), .B(n619), .C(n618), .Z(n511) );
  AO6SVTX8 U1323 ( .A(n1531), .B(n1508), .C(n506), .Z(n619) );
  ND2SVTX4 U1324 ( .A(n996), .B(n1114), .Z(n997) );
  ND4ABCSVTX8 U1325 ( .A(n1284), .B(n1283), .C(n1362), .D(n764), .Z(n805) );
  ND3ABSVTX8 U1326 ( .A(n1451), .B(n482), .C(n1398), .Z(n481) );
  IVSVTX4 U1327 ( .A(n1434), .Z(n482) );
  ND2SVTX4 U1328 ( .A(n350), .B(n1201), .Z(n485) );
  IVSVTX4 U1329 ( .A(n1109), .Z(n1104) );
  NR2SVTX8 U1330 ( .A(n358), .B(n1052), .Z(n486) );
  IVSVTX4 U1331 ( .A(n1052), .Z(n1276) );
  IVSVTX10 U1332 ( .A(n1143), .Z(n1172) );
  IVSVTX4 U1333 ( .A(n494), .Z(n1199) );
  NR3SVTX8 U1334 ( .A(n497), .B(n638), .C(n500), .Z(n825) );
  AO7SVTX8 U1335 ( .A(n499), .B(n1390), .C(n498), .Z(n500) );
  ND3SVTX8 U1336 ( .A(n350), .B(n1166), .C(n1167), .Z(n499) );
  ND2SVTX8 U1337 ( .A(n502), .B(n501), .Z(n1516) );
  ND2ASVTX6 U1338 ( .A(n230), .B(n1516), .Z(n1529) );
  NR2ASVTX8 U1339 ( .A(n230), .B(n1516), .Z(n1528) );
  ND2SVTX6 U1340 ( .A(n1519), .B(n1506), .Z(n1537) );
  ND3SVTX8 U1341 ( .A(n602), .B(n232), .C(n601), .Z(n505) );
  AO6SVTX6 U1342 ( .A(n506), .B(n1491), .C(n1490), .Z(n537) );
  AO7SVTX8 U1343 ( .A(n1536), .B(n539), .C(n538), .Z(n506) );
  AO6SVTX8 U1344 ( .A(n1236), .B(n231), .C(n509), .Z(n508) );
  ND2SVTX6 U1345 ( .A(n1102), .B(n1101), .Z(n1236) );
  ND3ABSVTX8 U1346 ( .A(n1149), .B(n998), .C(n997), .Z(n1041) );
  NR2SVTX8 U1347 ( .A(n513), .B(n1177), .Z(n904) );
  NR2SVTX4 U1348 ( .A(n941), .B(n682), .Z(n513) );
  ND2SVTX6 U1349 ( .A(n1071), .B(n850), .Z(n1219) );
  NR2SVTX8 U1350 ( .A(O[29]), .B(n904), .Z(n515) );
  IVSVTX4 U1351 ( .A(n1277), .Z(n516) );
  NR2ASVTX6 U1352 ( .A(n1196), .B(n1411), .Z(n1277) );
  NR2SVTX4 U1353 ( .A(n518), .B(n960), .Z(n1072) );
  ND2SVTX6 U1354 ( .A(n331), .B(n1355), .Z(n1470) );
  ND3SVTX6 U1355 ( .A(n1470), .B(n524), .C(n523), .Z(n1700) );
  ND2ASVTX8 U1356 ( .A(n1232), .B(n532), .Z(n534) );
  IVSVTX4 U1357 ( .A(n1231), .Z(n532) );
  ND2SVTX8 U1358 ( .A(n635), .B(n1230), .Z(n1231) );
  ND2SVTX8 U1359 ( .A(n673), .B(n533), .Z(n1230) );
  ND2SVTX8 U1360 ( .A(n535), .B(n1046), .Z(n1232) );
  ND2ASVTX8 U1361 ( .A(O[27]), .B(n672), .Z(n535) );
  ND2ASVTX8 U1362 ( .A(n358), .B(n542), .Z(n1046) );
  ND2SVTX6 U1363 ( .A(n537), .B(n536), .Z(n1489) );
  ND3SVTX8 U1364 ( .A(n1491), .B(n1508), .C(n1531), .Z(n536) );
  AO7SVTX8 U1365 ( .A(n1488), .B(n1653), .C(n1487), .Z(n1531) );
  ND4ABSVTX6 U1366 ( .A(n1726), .B(n1549), .C(n782), .D(n247), .Z(n1532) );
  ND2ASVTX6 U1367 ( .A(n289), .B(n1501), .Z(n1582) );
  ND2SVTX6 U1368 ( .A(n845), .B(n1533), .Z(n539) );
  ND2SVTX8 U1369 ( .A(n1205), .B(n1133), .Z(n541) );
  ND3SVTX8 U1370 ( .A(n635), .B(n634), .C(n1046), .Z(n1047) );
  ND3SVTX8 U1371 ( .A(n1043), .B(n1044), .C(n543), .Z(n542) );
  ND2SVTX8 U1372 ( .A(n891), .B(n1100), .Z(n1043) );
  ND2SVTX4 U1373 ( .A(n544), .B(n545), .Z(n1225) );
  IVSVTX4 U1374 ( .A(n724), .Z(n545) );
  ND2SVTX4 U1375 ( .A(n1280), .B(n1207), .Z(n544) );
  AO4SVTX6 U1376 ( .A(n889), .B(n1353), .C(n254), .D(n534), .Z(n547) );
  ND3SVTX8 U1377 ( .A(n1327), .B(n1326), .C(n1346), .Z(n1259) );
  AO4SVTX8 U1378 ( .A(n381), .B(n859), .C(n350), .D(n551), .Z(n1326) );
  ND2ASVTX8 U1379 ( .A(n552), .B(n1175), .Z(n1207) );
  ND2SVTX8 U1380 ( .A(n219), .B(n960), .Z(n1175) );
  ND2SVTX6 U1381 ( .A(n555), .B(n568), .Z(n554) );
  IVSVTX4 U1382 ( .A(n556), .Z(n566) );
  IVSVTX4 U1383 ( .A(n558), .Z(n564) );
  AO6CSVTX8 U1384 ( .A(n1382), .B(n248), .C(n560), .Z(n561) );
  AO7SVTX8 U1385 ( .A(n1381), .B(n1380), .C(n874), .Z(n562) );
  ND2SVTX6 U1386 ( .A(n570), .B(n566), .Z(n565) );
  IVSVTX4 U1387 ( .A(n1443), .Z(n570) );
  EO3SVTX8 U1388 ( .A(n573), .B(n572), .C(n581), .Z(n1587) );
  ND2SVTX6 U1389 ( .A(n1579), .B(n1580), .Z(n572) );
  ND2SVTX8 U1390 ( .A(n642), .B(n574), .Z(n1665) );
  NR2ASVTX6 U1391 ( .A(n1377), .B(n574), .Z(n1378) );
  ND2SVTX1 U1392 ( .A(n1498), .B(n575), .Z(n1494) );
  NR2SVTX8 U1393 ( .A(n1231), .B(n1232), .Z(n578) );
  EO3SVTX8 U1394 ( .A(n1527), .B(n633), .C(n590), .Z(n1594) );
  IVSVTX4 U1395 ( .A(n1503), .Z(n579) );
  NR2SVTX8 U1396 ( .A(n939), .B(n633), .Z(n581) );
  IVSVTX4 U1397 ( .A(n583), .Z(n681) );
  NR2SVTX6 U1398 ( .A(n1240), .B(n583), .Z(n678) );
  AO6CSVTX8 U1399 ( .A(n1372), .B(n1371), .C(n250), .Z(n1381) );
  ND2SVTX6 U1400 ( .A(n721), .B(n720), .Z(n1382) );
  AO7SVTX8 U1401 ( .A(n688), .B(n588), .C(n587), .Z(n1545) );
  ENSVTX8 U1402 ( .A(n230), .B(n589), .Z(n1250) );
  IVSVTX4 U1403 ( .A(n633), .Z(n592) );
  ND2SVTX4 U1404 ( .A(n592), .B(n1544), .Z(n632) );
  IVSVTX4 U1405 ( .A(n591), .Z(n1567) );
  NR2SVTX8 U1406 ( .A(n415), .B(n1052), .Z(n593) );
  ND2SVTX4 U1407 ( .A(n914), .B(n239), .Z(n617) );
  NR2SVTX8 U1408 ( .A(n1265), .B(n1437), .Z(n1311) );
  MUX21NSVTX8 U1409 ( .A(n1158), .B(n1164), .S(n1221), .Z(n1437) );
  MUX21NSVTX8 U1410 ( .A(n1127), .B(n1126), .S(n748), .Z(n1158) );
  ND2SVTX4 U1411 ( .A(n597), .B(n1309), .Z(n1265) );
  NR2SVTX4 U1412 ( .A(n1595), .B(n1594), .Z(n626) );
  ND2ASVTX8 U1413 ( .A(n511), .B(n1521), .Z(n633) );
  ND2SVTX4 U1414 ( .A(n1526), .B(n621), .Z(n599) );
  AO1SVTX6 U1415 ( .A(n742), .B(n1228), .C(n1443), .D(n648), .Z(n600) );
  NR2SVTX8 U1416 ( .A(n1519), .B(n1506), .Z(n1534) );
  EO3SVTX8 U1417 ( .A(n881), .B(n604), .C(n1585), .Z(n1588) );
  ND2SVTX8 U1418 ( .A(n605), .B(n1249), .Z(n855) );
  NR2SVTX8 U1419 ( .A(N[22]), .B(N[25]), .Z(n609) );
  NR3ABSVTX8 U1420 ( .A(n1315), .B(n1316), .C(n610), .Z(n1210) );
  NR3ABSVTX8 U1421 ( .A(n1342), .B(n1341), .C(n611), .Z(n1209) );
  ND2SVTX4 U1422 ( .A(n1205), .B(n1325), .Z(n1334) );
  ND2SVTX4 U1423 ( .A(n612), .B(n1203), .Z(n1341) );
  NR2SVTX4 U1424 ( .A(n814), .B(n1204), .Z(n612) );
  ND2ASVTX8 U1425 ( .A(n815), .B(n924), .Z(n1052) );
  AO7SVTX6 U1426 ( .A(n884), .B(n614), .C(n613), .Z(n1501) );
  F_ENSVTX2 U1427 ( .A(n675), .B(n831), .Z(n614) );
  IVSVTX4 U1428 ( .A(n1498), .Z(n1301) );
  ENSVTX4 U1429 ( .A(n1524), .B(n621), .Z(n1592) );
  IVSVTX4 U1430 ( .A(n1615), .Z(n1608) );
  ND2SVTX4 U1431 ( .A(n1592), .B(n1593), .Z(n630) );
  AO7SVTX6 U1432 ( .A(n1643), .B(n1569), .C(n1644), .Z(n1635) );
  ND2SVTX4 U1433 ( .A(n1568), .B(n628), .Z(n1644) );
  IVSVTX4 U1434 ( .A(n1571), .Z(n629) );
  IVSVTX4 U1435 ( .A(n632), .Z(n1568) );
  AO7SVTX8 U1436 ( .A(n521), .B(n1405), .C(n636), .Z(n1416) );
  ND2SVTX6 U1437 ( .A(n778), .B(n240), .Z(n1253) );
  ND2SVTX4 U1438 ( .A(n791), .B(n240), .Z(n779) );
  ND2SVTX4 U1439 ( .A(n706), .B(n705), .Z(n1288) );
  ND3ABSVTX8 U1440 ( .A(n1286), .B(n1285), .C(n640), .Z(n705) );
  AO7SVTX6 U1441 ( .A(n1285), .B(n855), .C(n1286), .Z(n706) );
  IVSVTX4 U1442 ( .A(n213), .Z(n1247) );
  ND4ABSVTX8 U1443 ( .A(n658), .B(n657), .C(n655), .D(n656), .Z(n856) );
  NR2SVTX6 U1444 ( .A(n1510), .B(n684), .Z(n645) );
  ND2SVTX6 U1445 ( .A(n646), .B(n647), .Z(n1462) );
  ND2SVTX8 U1446 ( .A(n232), .B(n1322), .Z(n647) );
  ND4ABSVTX8 U1447 ( .A(n1461), .B(n1321), .C(n1460), .D(n647), .Z(n1695) );
  AO7ABSVTX4 U1448 ( .A(n241), .B(n1270), .C(n1269), .Z(n1271) );
  IVSVTX4 U1449 ( .A(n1346), .Z(n1318) );
  IVSVTX4 U1450 ( .A(n1253), .Z(n1194) );
  ND2SVTX4 U1451 ( .A(n761), .B(n1305), .Z(n831) );
  IVSVTX8 U1452 ( .A(n1665), .Z(n1676) );
  IVSVTX10 U1453 ( .A(n1008), .Z(n989) );
  ND2SVTX4 U1454 ( .A(n650), .B(n649), .Z(n1497) );
  ND2SVTX2 U1455 ( .A(n249), .B(n1245), .Z(n1233) );
  ND2SVTX4 U1456 ( .A(n653), .B(n249), .Z(n652) );
  ND2SVTX4 U1457 ( .A(n231), .B(n783), .Z(n655) );
  NR2ASVTX6 U1458 ( .A(n1267), .B(n1184), .Z(n657) );
  NR2ASVTX6 U1459 ( .A(n1222), .B(n1109), .Z(n658) );
  AN3SVTX6 U1460 ( .A(n804), .B(n660), .C(n925), .Z(n654) );
  ND2SVTX6 U1461 ( .A(n967), .B(n966), .Z(n785) );
  AO7SVTX6 U1462 ( .A(n435), .B(n838), .C(n837), .Z(n672) );
  ND2ASVTX8 U1463 ( .A(n1137), .B(n1004), .Z(n1057) );
  AO7SVTX6 U1464 ( .A(n829), .B(n999), .C(n665), .Z(n778) );
  ND2SVTX4 U1465 ( .A(n942), .B(n475), .Z(n955) );
  ND3SVTX6 U1466 ( .A(n981), .B(n958), .C(n957), .Z(n956) );
  ND2SVTX4 U1467 ( .A(n1026), .B(n1030), .Z(n667) );
  ND2SVTX4 U1468 ( .A(n669), .B(n668), .Z(n1081) );
  AO2SVTX6 U1469 ( .A(n910), .B(n240), .C(n1093), .D(n891), .Z(n1078) );
  NR2SVTX4 U1470 ( .A(n1736), .B(n1455), .Z(n1457) );
  ND3ABSVTX8 U1471 ( .A(n888), .B(n1230), .C(n671), .Z(n1436) );
  IVSVTX10 U1472 ( .A(n674), .Z(n872) );
  ND2ASVTX8 U1473 ( .A(n1230), .B(n1047), .Z(n674) );
  ND2ASVTX8 U1474 ( .A(n743), .B(n742), .Z(n741) );
  ND2ASVTX8 U1475 ( .A(n977), .B(n683), .Z(n792) );
  AO2ABSVTX8 U1476 ( .C(n989), .D(n683), .A(n1172), .B(n1039), .Z(n690) );
  ND2SVTX4 U1477 ( .A(n240), .B(n1093), .Z(n692) );
  NR2SVTX4 U1478 ( .A(n234), .B(n724), .Z(n691) );
  ND2SVTX4 U1479 ( .A(n830), .B(n1094), .Z(n693) );
  ND2SVTX4 U1480 ( .A(n891), .B(n1214), .Z(n694) );
  ND3ABSVTX8 U1481 ( .A(n856), .B(n1293), .C(n1112), .Z(n695) );
  ND2SVTX6 U1482 ( .A(n1519), .B(n855), .Z(n699) );
  NR2SVTX6 U1483 ( .A(n697), .B(n855), .Z(n696) );
  AO8SVTX8 U1484 ( .A(n698), .B(n248), .C(n227), .D(n1287), .Z(n797) );
  ND2ASVTX8 U1485 ( .A(n1247), .B(n701), .Z(n703) );
  NR2SVTX4 U1486 ( .A(n805), .B(n710), .Z(n708) );
  IVSVTX4 U1487 ( .A(n815), .Z(n714) );
  ND2SVTX8 U1488 ( .A(n716), .B(n715), .Z(n1214) );
  IVSVTX4 U1489 ( .A(n814), .Z(n719) );
  AO21DSVTX8 U1490 ( .A(n1360), .B(n1369), .C(n722), .D(n1289), .Z(n721) );
  ND2SVTX4 U1491 ( .A(n725), .B(n540), .Z(n1315) );
  ND2SVTX4 U1492 ( .A(n1324), .B(n1345), .Z(n1211) );
  AN2SVTX8 U1493 ( .A(n714), .B(n1196), .Z(n1208) );
  NR2ASVTX6 U1494 ( .A(n1279), .B(n1186), .Z(n1212) );
  ND4ABSVTX8 U1495 ( .A(n1475), .B(n1476), .C(n726), .D(n1477), .Z(n1686) );
  AO7SVTX4 U1496 ( .A(n884), .B(n727), .C(n1304), .Z(n1499) );
  ND2SVTX4 U1497 ( .A(n640), .B(n742), .Z(n1302) );
  NR2SVTX4 U1498 ( .A(n1384), .B(n1386), .Z(n758) );
  NR2SVTX8 U1499 ( .A(n1401), .B(n1408), .Z(n1386) );
  ND3ABSVTX8 U1500 ( .A(n259), .B(n1135), .C(n358), .Z(n732) );
  NR2SVTX4 U1501 ( .A(n257), .B(n870), .Z(n1402) );
  IVSVTX4 U1502 ( .A(n1310), .Z(n1141) );
  NR2ASVTX6 U1503 ( .A(n1368), .B(n1369), .Z(n1372) );
  NR2ASVTX6 U1504 ( .A(n737), .B(n1597), .Z(n1602) );
  ND2SVTX6 U1505 ( .A(n738), .B(n739), .Z(n1504) );
  AO2SVTX2 U1506 ( .A(n1578), .B(n1546), .C(n496), .D(n448), .Z(n739) );
  ND3ABSVTX8 U1507 ( .A(n866), .B(n1229), .C(n1249), .Z(n743) );
  IVSVTX4 U1508 ( .A(n1275), .Z(n746) );
  IVSVTX4 U1509 ( .A(n1130), .Z(n1131) );
  ND2ASVTX8 U1510 ( .A(n1429), .B(n1459), .Z(n1697) );
  ENSVTX4 U1511 ( .A(n237), .B(n1369), .Z(n1322) );
  IVSVTX10 U1512 ( .A(n1443), .Z(n921) );
  NR2SVTX4 U1513 ( .A(n540), .B(n752), .Z(n1042) );
  AO7ASVTX8 U1514 ( .A(n1136), .B(n1408), .C(n1138), .Z(n1140) );
  BFSVTX6 U1515 ( .A(n1396), .Z(n754) );
  ND2SVTX4 U1516 ( .A(n1434), .B(n1398), .Z(n755) );
  NR2SVTX4 U1517 ( .A(n1449), .B(n754), .Z(n1434) );
  NR3ABSVTX8 U1518 ( .A(n759), .B(n758), .C(n757), .Z(n1394) );
  ND2SVTX6 U1519 ( .A(n1227), .B(n760), .Z(n756) );
  ND2SVTX8 U1520 ( .A(n742), .B(n740), .Z(n763) );
  ND2SVTX6 U1521 ( .A(n762), .B(n1244), .Z(n1246) );
  NR3SVTX6 U1522 ( .A(n326), .B(n765), .C(n766), .Z(n1283) );
  ENSVTX8 U1523 ( .A(n252), .B(n855), .Z(n767) );
  ND2SVTX6 U1524 ( .A(n769), .B(n768), .Z(n895) );
  NR2SVTX6 U1525 ( .A(N[25]), .B(N[26]), .Z(n768) );
  BFSVTX6 U1526 ( .A(n856), .Z(n770) );
  ND2SVTX4 U1527 ( .A(n770), .B(n1554), .Z(n1290) );
  AO5ASVTX8 U1528 ( .B(n877), .A(n252), .C(n1565), .Z(n771) );
  ND3SVTX6 U1529 ( .A(n959), .B(N[7]), .C(n960), .Z(n774) );
  ND2SVTX6 U1530 ( .A(n774), .B(n773), .Z(n1222) );
  IVSVTX2 U1531 ( .A(n1083), .Z(n773) );
  ND2SVTX4 U1532 ( .A(n1048), .B(n792), .Z(n791) );
  ND2SVTX4 U1533 ( .A(n830), .B(n914), .Z(n780) );
  AO2SVTX6 U1534 ( .A(n778), .B(n891), .C(n1099), .D(n1136), .Z(n781) );
  NR2SVTX4 U1535 ( .A(n1549), .B(n1291), .Z(n1308) );
  NR2ASVTX6 U1536 ( .A(n251), .B(n839), .Z(n1549) );
  ND2SVTX6 U1537 ( .A(n798), .B(n797), .Z(n1554) );
  ND2SVTX6 U1538 ( .A(n847), .B(n848), .Z(n1307) );
  ND2SVTX4 U1539 ( .A(n840), .B(n839), .Z(n1660) );
  NR2SVTX4 U1540 ( .A(n1247), .B(n875), .Z(n784) );
  ND2SVTX4 U1541 ( .A(n1280), .B(n785), .Z(n968) );
  NR2ASVTX6 U1542 ( .A(N[3]), .B(n786), .Z(n1050) );
  ND2ASVTX8 U1543 ( .A(n1084), .B(n960), .Z(n786) );
  ENSVTX8 U1544 ( .A(n255), .B(n787), .Z(n1441) );
  IVSVTX6 U1545 ( .A(N[14]), .Z(n1008) );
  NR2ASVTX6 U1546 ( .A(n256), .B(n1418), .Z(n789) );
  BFSVTX6 U1547 ( .A(n789), .Z(n790) );
  IVSVTX4 U1548 ( .A(n899), .Z(n900) );
  ND2SVTX6 U1549 ( .A(n795), .B(n794), .Z(n992) );
  NR2SVTX6 U1550 ( .A(N[9]), .B(N[10]), .Z(n795) );
  ND2SVTX6 U1551 ( .A(n264), .B(n945), .Z(n1067) );
  NR2SVTX4 U1552 ( .A(n358), .B(n799), .Z(n1181) );
  IVSVTX4 U1553 ( .A(n800), .Z(n1149) );
  IVSVTX4 U1554 ( .A(n1286), .Z(n801) );
  ND2SVTX6 U1555 ( .A(n1219), .B(n239), .Z(n803) );
  NR2ASVTX8 U1556 ( .A(n253), .B(n1573), .Z(n1296) );
  ND2SVTX8 U1557 ( .A(n809), .B(n808), .Z(n1573) );
  ND2SVTX8 U1558 ( .A(n232), .B(n1250), .Z(n808) );
  ND2SVTX4 U1559 ( .A(n811), .B(n812), .Z(n943) );
  NR2SVTX4 U1560 ( .A(N[13]), .B(N[15]), .Z(n811) );
  NR2SVTX4 U1561 ( .A(N[12]), .B(N[14]), .Z(n812) );
  ND2SVTX8 U1562 ( .A(n816), .B(n817), .Z(n1763) );
  IVSVTX4 U1563 ( .A(n822), .Z(n1174) );
  ND2SVTX4 U1564 ( .A(n1280), .B(n822), .Z(n819) );
  IVSVTX6 U1565 ( .A(n946), .Z(n1117) );
  ND2SVTX4 U1566 ( .A(n245), .B(n666), .Z(n827) );
  ND2SVTX8 U1567 ( .A(n828), .B(n453), .Z(n947) );
  AO20SVTX8 U1568 ( .A(n1381), .B(n1380), .C(n921), .D(n1374), .Z(n1375) );
  ND2ASVTX8 U1569 ( .A(n478), .B(n1435), .Z(n833) );
  ND2SVTX4 U1570 ( .A(n232), .B(n1442), .Z(n834) );
  NR2SVTX8 U1571 ( .A(n1107), .B(n1186), .Z(n1258) );
  ND2SVTX8 U1572 ( .A(n1090), .B(n934), .Z(n1213) );
  ND2SVTX6 U1573 ( .A(n1357), .B(n1356), .Z(n841) );
  IVSVTX4 U1574 ( .A(n841), .Z(n1358) );
  IVSVTX4 U1575 ( .A(n846), .Z(n1228) );
  IVSVTX4 U1576 ( .A(n1268), .Z(n1270) );
  NR2SVTX4 U1577 ( .A(N[30]), .B(N[28]), .Z(n851) );
  ND2SVTX6 U1578 ( .A(n1700), .B(n1702), .Z(n1474) );
  ND2SVTX6 U1579 ( .A(n860), .B(n861), .Z(n1252) );
  ND4SVTX6 U1580 ( .A(n1366), .B(n1363), .C(n1364), .D(n1365), .Z(n1370) );
  BFSVTX2 U1581 ( .A(n1667), .Z(n864) );
  IVSVTX4 U1582 ( .A(n1267), .Z(n1191) );
  ND2ASVTX8 U1583 ( .A(n1199), .B(n1200), .Z(n1267) );
  AO7SVTX4 U1584 ( .A(n1019), .B(n1020), .C(n1114), .Z(n1028) );
  MUX21NSVTX8 U1585 ( .A(n882), .B(n865), .S(n748), .Z(n1132) );
  ND3ASVTX4 U1586 ( .A(N[10]), .B(n977), .C(n1005), .Z(n948) );
  BFSVTX2 U1587 ( .A(n1437), .Z(n1451) );
  IVSVTX0H U1588 ( .A(n1678), .Z(n868) );
  AN4SVTX8 U1589 ( .A(n814), .B(n879), .C(n870), .D(n1207), .Z(n878) );
  NR3ASVTX6 U1590 ( .A(n1345), .B(n1340), .C(n1338), .Z(n1323) );
  NR2ASVTX4 U1591 ( .A(n398), .B(n815), .Z(n1049) );
  ND2ASVTX8 U1592 ( .A(n1480), .B(n1383), .Z(n919) );
  CTIVSVTX2 U1593 ( .A(n870), .Z(n1147) );
  ND3ASVTX4 U1594 ( .A(n1029), .B(n1010), .C(n1009), .Z(n1012) );
  IVSVTX2 U1595 ( .A(n438), .Z(n1029) );
  AO7SVTX2 U1596 ( .A(n1087), .B(n1084), .C(n475), .Z(n1003) );
  F_IVSVTX1 U1597 ( .A(n1750), .Z(n1759) );
  EOSVTX2 U1598 ( .A(n1583), .B(n619), .Z(n883) );
  F_ND2SVTX0H U1599 ( .A(n1088), .B(n1143), .Z(n1089) );
  MUX21NSVTX2 U1600 ( .A(n1236), .B(n1235), .S(n231), .Z(n1237) );
  AO2SVTX4 U1601 ( .A(n791), .B(n830), .C(n891), .D(n914), .Z(n1102) );
  FAS1SVTX2 U1602 ( .A(n1575), .B(n1574), .CI(n463), .CO(n1517), .Z(n1584) );
  OR2SVTX4 U1603 ( .A(n1231), .B(n1232), .Z(n886) );
  ND3ABSVTX4 U1604 ( .A(n1402), .B(n867), .C(n932), .Z(n1419) );
  IVSVTX4 U1605 ( .A(n1117), .Z(n890) );
  IVSVTX12 U1606 ( .A(n872), .Z(n1248) );
  ND2SVTX4 U1607 ( .A(n424), .B(n1318), .Z(n1319) );
  ND2SVTX6 U1608 ( .A(n264), .B(n945), .Z(n893) );
  NR3SVTX6 U1609 ( .A(n438), .B(n245), .C(n949), .Z(n950) );
  IVSVTX4 U1610 ( .A(n1627), .Z(n906) );
  ND2SVTX4 U1611 ( .A(n873), .B(n496), .Z(n1503) );
  ND2ASVTX8 U1612 ( .A(n1148), .B(n1147), .Z(n1309) );
  IVSVTX2 U1613 ( .A(n1261), .Z(n1263) );
  ND2SVTX4 U1614 ( .A(n995), .B(n994), .Z(n996) );
  IVSVTX2 U1615 ( .A(n1219), .Z(n1108) );
  F_ND2ASVTX2 U1616 ( .A(n1135), .B(n1145), .Z(n1120) );
  NR3SVTX6 U1617 ( .A(n1180), .B(n1165), .C(n1163), .Z(n1261) );
  B_ND2SVTX0H U1618 ( .A(N[2]), .B(n422), .Z(n1173) );
  IVSVTX4 U1619 ( .A(n1574), .Z(n1286) );
  ND2SVTX2 U1620 ( .A(n1280), .B(n1279), .Z(n1281) );
  AO6SVTX1 U1621 ( .A(n1540), .B(n1560), .C(n1539), .Z(n1541) );
  IVSVTX2 U1622 ( .A(N[19]), .Z(n942) );
  IVSVTX2 U1623 ( .A(n1710), .Z(n1704) );
  AO7SVTX2 U1624 ( .A(n1009), .B(n959), .C(n437), .Z(n964) );
  AO7SVTX2 U1625 ( .A(n262), .B(n990), .C(n1146), .Z(n993) );
  NR2ASVTX2 U1626 ( .A(N[0]), .B(n959), .Z(n1086) );
  IVSVTX2 U1627 ( .A(n1061), .Z(n1062) );
  IVSVTX2 U1628 ( .A(n1233), .Z(n1234) );
  ND2SVTX2 U1629 ( .A(n1251), .B(n1332), .Z(n1328) );
  IVSVTX4 U1630 ( .A(n496), .Z(n1513) );
  IVSVTX2 U1631 ( .A(n1480), .Z(n1481) );
  F_ND2SVTX0H U1632 ( .A(n1735), .B(n1734), .Z(n1738) );
  F_ND2SVTX1 U1633 ( .A(n1454), .B(n1716), .Z(n1725) );
  ND4ABSVTX4 U1634 ( .A(n521), .B(n675), .C(n1303), .D(n1305), .Z(n1304) );
  ND2SVTX4 U1635 ( .A(n830), .B(n1093), .Z(n1066) );
  AO7SVTX1 U1636 ( .A(n1538), .B(n445), .C(n1537), .Z(n1539) );
  IVSVTX4 U1637 ( .A(n1176), .Z(n1116) );
  ND2SVTX4 U1638 ( .A(n1214), .B(n830), .Z(n1092) );
  F_ND2SVTX1 U1639 ( .A(n1740), .B(n1739), .Z(n1743) );
  NR2SVTX2 U1640 ( .A(n1172), .B(n1054), .Z(n1055) );
  ND2SVTX4 U1641 ( .A(n873), .B(n1435), .Z(n1430) );
  F_ND2SVTX1 U1642 ( .A(n1685), .B(n461), .Z(n1694) );
  AN2SVTX4 U1643 ( .A(n1613), .B(n1614), .Z(n1610) );
  IVSVTX4 U1644 ( .A(n1552), .Z(n899) );
  BFSVTX2 U1645 ( .A(n1639), .Z(n901) );
  F_AN2SVTX2 U1646 ( .A(n1280), .B(n1207), .Z(n903) );
  AO3SVTX2 U1647 ( .A(n431), .B(n1221), .C(n597), .D(n1309), .Z(n1458) );
  AO7ASVTX4 U1648 ( .A(n1049), .B(n791), .C(n1221), .Z(n1051) );
  AO7ABSVTX8 U1649 ( .A(n1251), .B(n1275), .C(n1274), .Z(n1368) );
  AO7NSVTX4 U1650 ( .A(n1423), .B(n1750), .C(n1422), .Z(n923) );
  ND2SVTX4 U1651 ( .A(n906), .B(n907), .Z(n909) );
  ND2SVTX4 U1652 ( .A(n908), .B(n909), .Z(O[25]) );
  AO7SVTX8 U1653 ( .A(n1463), .B(n1462), .C(n1461), .Z(n1696) );
  ND2SVTX2 U1654 ( .A(n967), .B(n966), .Z(n910) );
  ND2SVTX2 U1655 ( .A(n766), .B(n1220), .Z(n1269) );
  AO7ABSVTX4 U1656 ( .A(n424), .B(n1329), .C(n1328), .Z(n1349) );
  AO6SVTX8 U1657 ( .A(n1667), .B(n1486), .C(n1485), .Z(n1487) );
  AO7SVTX8 U1658 ( .A(n1464), .B(n1697), .C(n1696), .Z(n1465) );
  IVSVTX2 U1659 ( .A(n1449), .Z(n1400) );
  ENSVTX4 U1660 ( .A(n913), .B(n1646), .Z(O[18]) );
  AO6CSVTX8 U1661 ( .A(n1631), .B(n1616), .C(n1608), .Z(n1617) );
  AO6CSVTX8 U1662 ( .A(n1631), .B(n451), .C(n915), .Z(n1622) );
  AO6SVTX1 U1663 ( .A(n1560), .B(n1559), .C(n449), .Z(n1561) );
  AO7SVTX8 U1664 ( .A(n1297), .B(n1296), .C(n1295), .Z(n1558) );
  ND2ASVTX8 U1665 ( .A(n246), .B(n1627), .Z(n1628) );
  ENSVTX8 U1666 ( .A(n228), .B(n1622), .Z(O[22]) );
  ND2SVTX2 U1667 ( .A(n682), .B(n1036), .Z(n917) );
  NR2ASVTX4 U1668 ( .A(n1151), .B(n682), .Z(n1070) );
  BFSVTX2 U1669 ( .A(n682), .Z(O[30]) );
  AO1ABSVTX4 U1670 ( .A(n1039), .B(n999), .C(n963), .D(n962), .Z(n969) );
  ND2ASVTX4 U1671 ( .A(n1400), .B(n1450), .Z(n1735) );
  AO7SVTX1 U1672 ( .A(n884), .B(n623), .C(n875), .Z(n1624) );
  ND2SVTX4 U1673 ( .A(n1327), .B(n1326), .Z(n1332) );
  NR2SVTX2 U1674 ( .A(n1172), .B(n1058), .Z(n1060) );
  NR2ASVTX6 U1675 ( .A(N[8]), .B(n1172), .Z(n1176) );
  ND2SVTX4 U1676 ( .A(N[7]), .B(n973), .Z(n974) );
  ND2SVTX4 U1677 ( .A(n920), .B(n1521), .Z(n1548) );
  F_IVSVTX0H U1678 ( .A(n1618), .Z(n1619) );
  AO7SVTX4 U1679 ( .A(n496), .B(n1578), .C(n684), .Z(n1579) );
  F_MUX21NSVTX1 U1680 ( .A(n873), .B(n1510), .S(n1578), .Z(n1492) );
  ND2SVTX2 U1681 ( .A(n1520), .B(n1578), .Z(n1523) );
  ND2SVTX4 U1682 ( .A(n403), .B(n426), .Z(n1395) );
  OR2SVTX4 U1683 ( .A(n682), .B(n941), .Z(n927) );
  ND2SVTX4 U1684 ( .A(n1178), .B(n1084), .Z(n941) );
  AO6SVTX2 U1685 ( .A(n494), .B(n1200), .C(n1280), .Z(n1201) );
  ND2SVTX2 U1686 ( .A(n1243), .B(n740), .Z(n1244) );
  ND2SVTX4 U1687 ( .A(n1316), .B(n1315), .Z(n1338) );
  ENSVTX8 U1688 ( .A(n936), .B(n1611), .Z(O[24]) );
  ENSVTX8 U1689 ( .A(n938), .B(n1617), .Z(O[23]) );
  ND2SVTX2 U1690 ( .A(n1640), .B(n901), .Z(n1641) );
  NR2ASVTX1 U1691 ( .A(N[15]), .B(n1172), .Z(n1083) );
  F_ND2SVTX0H U1692 ( .A(N[18]), .B(n1143), .Z(n1073) );
  ENSVTX8 U1693 ( .A(n1629), .B(n1628), .Z(O[26]) );
  NR2ASVTX6 U1694 ( .A(n814), .B(n1198), .Z(n1163) );
  NR2ASVTX6 U1695 ( .A(N[7]), .B(n1159), .Z(n1198) );
  IVSVTX4 U1696 ( .A(n1145), .Z(n1159) );
  F_ND2SVTX1 U1697 ( .A(n1696), .B(n214), .Z(n1699) );
  IVSVTX0H U1698 ( .A(n1638), .Z(n1640) );
  ND3SVTX2 U1699 ( .A(n1342), .B(n1341), .C(n1317), .Z(n1344) );
  ND2SVTX2 U1700 ( .A(n1039), .B(N[19]), .Z(n970) );
  EOSVTX8 U1701 ( .A(n1505), .B(n1504), .Z(n1596) );
  BFSVTX2 U1702 ( .A(N[10]), .Z(n1142) );
  IVSVTX2 U1703 ( .A(n1531), .Z(n1552) );
  IVSVTX0H U1704 ( .A(N[8]), .Z(n1087) );
  F_AN2SVTX2 U1705 ( .A(n1613), .B(n1607), .Z(n938) );
  F_EOSVTX2 U1706 ( .A(n1564), .B(n1563), .Z(n940) );
  NR2ASVTX1 U1707 ( .A(N[0]), .B(n1172), .Z(n1139) );
  IVSVTX4 U1708 ( .A(N[17]), .Z(n981) );
  IVSVTX4 U1709 ( .A(N[25]), .Z(n1030) );
  IVSVTX4 U1710 ( .A(N[18]), .Z(n1026) );
  BFSVTX6 U1711 ( .A(N[6]), .Z(n1085) );
  IVSVTX4 U1712 ( .A(N[4]), .Z(n1115) );
  IVSVTX6 U1713 ( .A(N[5]), .Z(n1053) );
  NR2SVTX6 U1714 ( .A(n1067), .B(n947), .Z(n946) );
  IVSVTX4 U1715 ( .A(N[15]), .Z(n977) );
  IVSVTX4 U1716 ( .A(n948), .Z(n951) );
  NR2SVTX4 U1717 ( .A(N[23]), .B(N[21]), .Z(n953) );
  NR3SVTX8 U1718 ( .A(N[20]), .B(N[18]), .C(N[30]), .Z(n952) );
  IVSVTX4 U1719 ( .A(n1142), .Z(n1009) );
  ND3SVTX6 U1720 ( .A(n1146), .B(n1115), .C(n1053), .Z(n1014) );
  NR3SVTX8 U1721 ( .A(N[14]), .B(N[13]), .C(N[12]), .Z(n973) );
  ND2SVTX4 U1722 ( .A(n245), .B(n263), .Z(n978) );
  AO7SVTX4 U1723 ( .A(n979), .B(n978), .C(n977), .Z(n984) );
  ND3SVTX8 U1724 ( .A(n981), .B(n1023), .C(n980), .Z(n982) );
  NR3SVTX8 U1725 ( .A(n1000), .B(n1021), .C(n982), .Z(n983) );
  BFSVTX2 U1726 ( .A(N[26]), .Z(n987) );
  NR2SVTX6 U1727 ( .A(n992), .B(n991), .Z(n1016) );
  AO7SVTX1 U1728 ( .A(n1005), .B(n1084), .C(n453), .Z(n1007) );
  F_ND2SVTX0H U1729 ( .A(N[13]), .B(n1008), .Z(n1013) );
  ND3SVTX4 U1730 ( .A(n1013), .B(n1012), .C(n1011), .Z(n1020) );
  IVSVTX2 U1731 ( .A(n1014), .Z(n1015) );
  ND3SVTX2 U1732 ( .A(N[1]), .B(n262), .C(n1015), .Z(n1018) );
  NR2SVTX2 U1733 ( .A(n1018), .B(n1017), .Z(n1019) );
  ND2SVTX2 U1734 ( .A(N[21]), .B(n1039), .Z(n1025) );
  BFSVTX6 U1735 ( .A(N[17]), .Z(n1068) );
  IVSVTX2 U1736 ( .A(n1029), .Z(n1151) );
  ND2SVTX2 U1737 ( .A(n469), .B(n960), .Z(n1035) );
  ND2SVTX4 U1738 ( .A(n1085), .B(n1038), .Z(n1040) );
  IVSVTX4 U1739 ( .A(n1070), .Z(n1071) );
  NR2ASVTX2 U1740 ( .A(n914), .B(n1109), .Z(n1076) );
  NR2SVTX4 U1741 ( .A(n1076), .B(n1075), .Z(n1082) );
  NR2SVTX4 U1742 ( .A(n1109), .B(n302), .Z(n1098) );
  NR2SVTX4 U1743 ( .A(n242), .B(n1184), .Z(n1097) );
  ND4ABSVTX8 U1744 ( .A(n1097), .B(n1098), .C(n1095), .D(n1096), .Z(n1293) );
  NR2SVTX2 U1745 ( .A(n1235), .B(n826), .Z(n1111) );
  BFSVTX12 U1746 ( .A(n1117), .Z(n1154) );
  ND2ASVTX8 U1747 ( .A(n1106), .B(n1105), .Z(n1238) );
  ND2SVTX4 U1748 ( .A(n1120), .B(n1119), .Z(n1126) );
  ND2SVTX2 U1749 ( .A(N[5]), .B(n1154), .Z(n1122) );
  ND2SVTX4 U1750 ( .A(n1124), .B(n1123), .Z(n1388) );
  NR2SVTX8 U1751 ( .A(n1128), .B(n1396), .Z(n1310) );
  F_ND2ASVTX2 U1752 ( .A(n1137), .B(n1136), .Z(n1138) );
  NR3SVTX6 U1753 ( .A(n1198), .B(n1161), .C(n1160), .Z(n1165) );
  NR2SVTX4 U1754 ( .A(n1171), .B(n1174), .Z(n1169) );
  IVSVTX4 U1755 ( .A(n1217), .Z(n1190) );
  NR2ASVTX6 U1756 ( .A(n1216), .B(n1190), .Z(n1278) );
  ND2ASVTX8 U1757 ( .A(n1206), .B(n350), .Z(n1345) );
  ND2SVTX4 U1758 ( .A(n289), .B(n603), .Z(n1240) );
  ND2SVTX2 U1759 ( .A(n1299), .B(n249), .Z(n1241) );
  ND2SVTX4 U1760 ( .A(n428), .B(n1268), .Z(n1255) );
  ND2SVTX4 U1761 ( .A(n1256), .B(n1255), .Z(n1257) );
  NR2SVTX2 U1762 ( .A(n1278), .B(n1411), .Z(n1266) );
  ND2ASVTX8 U1763 ( .A(n1251), .B(n1273), .Z(n1274) );
  IVSVTX4 U1764 ( .A(n1278), .Z(n1279) );
  ND2ASVTX4 U1765 ( .A(n306), .B(n1307), .Z(n1728) );
  ND2ASVTX8 U1766 ( .A(n1247), .B(n1545), .Z(n1297) );
  ND2SVTX4 U1767 ( .A(n1294), .B(n1573), .Z(n1295) );
  IVSVTX4 U1768 ( .A(n1302), .Z(n1303) );
  IVSVTX4 U1769 ( .A(n1459), .Z(n1320) );
  ND2ASVTX8 U1770 ( .A(n1458), .B(n1320), .Z(n1731) );
  ND2SVTX4 U1771 ( .A(n1731), .B(n214), .Z(n1711) );
  ND2ASVTX8 U1772 ( .A(n1331), .B(n249), .Z(n1469) );
  NR2SVTX4 U1773 ( .A(n1336), .B(n1337), .Z(n1350) );
  NR2SVTX4 U1774 ( .A(n1711), .B(n1474), .Z(n1666) );
  ND2ASVTX8 U1775 ( .A(n1362), .B(n1368), .Z(n1480) );
  ND2SVTX4 U1776 ( .A(n921), .B(n1359), .Z(n1357) );
  ND2SVTX6 U1777 ( .A(n1652), .B(n461), .Z(n1673) );
  NR2SVTX4 U1778 ( .A(n1362), .B(n1361), .Z(n1366) );
  NR2SVTX4 U1779 ( .A(n1370), .B(n1369), .Z(n1367) );
  IVSVTX4 U1780 ( .A(n1370), .Z(n1371) );
  NR2SVTX8 U1781 ( .A(n1673), .B(n1484), .Z(n1486) );
  ND2SVTX4 U1782 ( .A(n1486), .B(n1666), .Z(n1488) );
  ND2SVTX4 U1783 ( .A(n1385), .B(n1387), .Z(n1417) );
  NR2SVTX2 U1784 ( .A(n259), .B(n1408), .Z(n1413) );
  AN2SVTX4 U1785 ( .A(n254), .B(n873), .Z(n1409) );
  NR3ABSVTX2 U1786 ( .A(N[0]), .B(n428), .C(n259), .Z(n1412) );
  AO6SVTX8 U1787 ( .A(n1414), .B(n1415), .C(n217), .Z(n1750) );
  ND2SVTX4 U1788 ( .A(n1417), .B(n1416), .Z(n1751) );
  IVSVTX4 U1789 ( .A(n1751), .Z(n1757) );
  AO7SVTX8 U1790 ( .A(n1423), .B(n1750), .C(n1422), .Z(n1717) );
  ND2ASVTX8 U1791 ( .A(n1399), .B(n1448), .Z(n1739) );
  AO6SVTX8 U1792 ( .A(n1717), .B(n1457), .C(n1456), .Z(n1653) );
  IVSVTX4 U1793 ( .A(n1695), .Z(n1464) );
  IVSVTX4 U1794 ( .A(n1460), .Z(n1463) );
  AO6SVTX8 U1795 ( .A(n919), .B(n1676), .C(n1482), .Z(n1483) );
  AO7SVTX8 U1796 ( .A(n1675), .B(n1484), .C(n1483), .Z(n1485) );
  ENSVTX8 U1797 ( .A(n1301), .B(n1489), .Z(n1578) );
  IVSVTX2 U1798 ( .A(n1623), .Z(n1496) );
  NR2SVTX4 U1799 ( .A(n1602), .B(n1605), .Z(n1599) );
  BFSVTX1 U1800 ( .A(n1506), .Z(n1518) );
  FAS1SVTX4 U1801 ( .A(n1519), .B(n1518), .CI(n1517), .CO(n1525), .Z(n1586) );
  F_ENSVTX2 U1802 ( .A(n1526), .B(n1525), .Z(n1524) );
  NR2SVTX4 U1803 ( .A(n1593), .B(n1592), .Z(n1620) );
  NR2SVTX4 U1804 ( .A(n1594), .B(n1595), .Z(n1618) );
  ND2SVTX4 U1805 ( .A(n1599), .B(n1614), .Z(n1601) );
  IVSVTX0H U1806 ( .A(n1536), .Z(n1560) );
  AO7SVTX2 U1807 ( .A(n1562), .B(n900), .C(n1561), .Z(n1563) );
  NR2SVTX8 U1808 ( .A(n1589), .B(n1588), .Z(n1632) );
  NR2SVTX4 U1809 ( .A(n1632), .B(n1638), .Z(n1591) );
  ND2SVTX4 U1810 ( .A(n1589), .B(n1588), .Z(n1633) );
  AO6SVTX8 U1811 ( .A(n1591), .B(n1635), .C(n1590), .Z(n1606) );
  ND2SVTX4 U1812 ( .A(n926), .B(n1596), .Z(n1607) );
  IVSVTX2 U1813 ( .A(n1602), .Z(n1603) );
  AO6SVTX8 U1814 ( .A(n1631), .B(n1610), .C(n1609), .Z(n1611) );
  ND2SVTX2 U1815 ( .A(n1624), .B(n1623), .Z(n1625) );
  IVSVTX2 U1816 ( .A(n1632), .Z(n1634) );
  ENSVTX4 U1817 ( .A(n1637), .B(n1636), .Z(O[20]) );
  EOSVTX4 U1818 ( .A(n1642), .B(n1641), .Z(O[19]) );
  IVSVTX0H U1819 ( .A(n1643), .Z(n1645) );
  ND2SVTX2 U1820 ( .A(n1645), .B(n1644), .Z(n1646) );
  IVSVTX2 U1821 ( .A(n1647), .Z(n1648) );
  ENSVTX4 U1822 ( .A(n1651), .B(n1650), .Z(O[17]) );
  BFSVTX1 U1823 ( .A(n1653), .Z(n1654) );
  IVSVTX4 U1824 ( .A(n1654), .Z(n1732) );
  EOSVTX4 U1825 ( .A(n1656), .B(n1655), .Z(O[10]) );
  AO7SVTX2 U1826 ( .A(n900), .B(n1726), .C(n1728), .Z(n1658) );
  ENSVTX4 U1827 ( .A(n1659), .B(n1658), .Z(O[15]) );
  ENSVTX4 U1828 ( .A(n1663), .B(n1662), .Z(O[16]) );
  ND2SVTX2 U1829 ( .A(n1677), .B(n1665), .Z(n1671) );
  IVSVTX2 U1830 ( .A(n1666), .Z(n1687) );
  IVSVTX2 U1831 ( .A(n864), .Z(n1689) );
  AO7SVTX1 U1832 ( .A(n902), .B(n1689), .C(n868), .Z(n1668) );
  AO6SVTX2 U1833 ( .A(n1669), .B(n1732), .C(n1668), .Z(n1670) );
  EOSVTX4 U1834 ( .A(n1671), .B(n1670), .Z(O[12]) );
  F_ND2SVTX1 U1835 ( .A(n919), .B(n1672), .Z(n1684) );
  IVSVTX2 U1836 ( .A(n1673), .Z(n1674) );
  NR2SVTX2 U1837 ( .A(n1687), .B(n1680), .Z(n1682) );
  IVSVTX0H U1838 ( .A(n1675), .Z(n1678) );
  AO6SVTX1 U1839 ( .A(n1678), .B(n1677), .C(n1676), .Z(n1679) );
  AO7SVTX1 U1840 ( .A(n1689), .B(n1680), .C(n1679), .Z(n1681) );
  AO6SVTX2 U1841 ( .A(n1682), .B(n1732), .C(n1681), .Z(n1683) );
  EOSVTX4 U1842 ( .A(n1684), .B(n1683), .Z(O[13]) );
  NR2SVTX2 U1843 ( .A(n1690), .B(n1687), .Z(n1692) );
  AO6SVTX2 U1844 ( .A(n1692), .B(n1732), .C(n1691), .Z(n1693) );
  EOSVTX4 U1845 ( .A(n1694), .B(n1693), .Z(O[11]) );
  AO6SVTX2 U1846 ( .A(n1732), .B(n412), .C(n1730), .Z(n1698) );
  EOSVTX4 U1847 ( .A(n1699), .B(n1698), .Z(O[7]) );
  NR2SVTX2 U1848 ( .A(n1704), .B(n1711), .Z(n1706) );
  AO6SVTX2 U1849 ( .A(n1732), .B(n1706), .C(n1705), .Z(n1707) );
  EOSVTX4 U1850 ( .A(n1708), .B(n1707), .Z(O[9]) );
  AO6SVTX2 U1851 ( .A(n1732), .B(n1713), .C(n1712), .Z(n1714) );
  EOSVTX4 U1852 ( .A(n1715), .B(n1714), .Z(O[8]) );
  IVSVTX1 U1853 ( .A(n310), .Z(n1718) );
  IVSVTX1 U1854 ( .A(n442), .Z(n1721) );
  AO6SVTX1 U1855 ( .A(n1721), .B(n1734), .C(n1720), .Z(n1722) );
  AO7SVTX2 U1856 ( .A(n923), .B(n1723), .C(n1722), .Z(n1724) );
  ENSVTX4 U1857 ( .A(n1725), .B(n1724), .Z(O[5]) );
  EOSVTX4 U1858 ( .A(n1729), .B(n900), .Z(O[14]) );
  ENSVTX4 U1859 ( .A(n1733), .B(n1732), .Z(O[6]) );
  AO7SVTX2 U1860 ( .A(n923), .B(n310), .C(n442), .Z(n1737) );
  AO7SVTX2 U1861 ( .A(n923), .B(n1741), .C(n443), .Z(n1742) );
  AO6SVTX2 U1862 ( .A(n1753), .B(n1759), .C(n1752), .Z(n1754) );
  EOSVTX4 U1863 ( .A(n1755), .B(n1754), .Z(O[1]) );
endmodule

