
module remap ( m1, m2 );
  input [27:0] m1;
  output [26:0] m2;
  wire   n1, n3, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n154, n155, n156, n157, n158, n160, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080;

  IVSVTX0H U3 ( .A(n1747), .Z(n1767) );
  AO6SVTX1 U4 ( .A(n2002), .B(n2036), .C(n596), .Z(n2031) );
  AO6SVTX1 U5 ( .A(n1992), .B(n174), .C(n22), .Z(n177) );
  AO2SVTX1 U6 ( .A(n2035), .B(n2036), .C(n599), .D(n528), .Z(n2075) );
  ENSVTX1 U7 ( .A(n1860), .B(n1859), .Z(n1895) );
  OR2SVTX2 U8 ( .A(n136), .B(n772), .Z(n815) );
  ND3SVTX4 U9 ( .A(n502), .B(n1920), .C(n663), .Z(n6) );
  EOSVTX0H U10 ( .A(n1718), .B(n219), .Z(n810) );
  EOSVTX0H U11 ( .A(n1434), .B(n1433), .Z(n1473) );
  AO6CSVTX2 U12 ( .A(n1670), .B(n1669), .C(n1668), .Z(n813) );
  AO6SVTX1 U13 ( .A(n1713), .B(n2036), .C(n597), .Z(n1714) );
  NR2ASVTX1 U14 ( .A(n1852), .B(n1851), .Z(n1860) );
  IVSVTX2 U15 ( .A(n1539), .Z(n336) );
  IVSVTX0H U16 ( .A(n1538), .Z(n1540) );
  EOSVTX1 U17 ( .A(n2042), .B(n2041), .Z(n2043) );
  ND3SVTX4 U18 ( .A(n1552), .B(n624), .C(n455), .Z(n623) );
  ND2SVTX2 U19 ( .A(n1922), .B(n1577), .Z(n1576) );
  ND3SVTX4 U20 ( .A(n1552), .B(n455), .C(n54), .Z(n626) );
  NR2ASVTX1 U21 ( .A(n299), .B(n44), .Z(n596) );
  ENSVTX0H U22 ( .A(n1773), .B(n1842), .Z(n1774) );
  EOSVTX0H U23 ( .A(n1381), .B(n1380), .Z(n1411) );
  EOSVTX1 U24 ( .A(n2021), .B(n2020), .Z(n2022) );
  EOSVTX0H U25 ( .A(n1439), .B(n1438), .Z(n1471) );
  ENSVTX0H U26 ( .A(n1369), .B(n1985), .Z(n772) );
  ND2ASVTX6 U27 ( .A(n635), .B(n587), .Z(n640) );
  ND2ASVTX6 U28 ( .A(n1426), .B(n286), .Z(n1915) );
  NR2ASVTX1 U29 ( .A(n2063), .B(n2062), .Z(n2068) );
  NR2ASVTX1 U30 ( .A(n1838), .B(n1837), .Z(n1844) );
  BFSVTX8 U31 ( .A(n1919), .Z(n223) );
  AO2SVTX1 U32 ( .A(n1467), .B(n1640), .C(n12), .D(n599), .Z(n1468) );
  NR2ASVTX1 U33 ( .A(n2045), .B(n2044), .Z(n2047) );
  AO6SVTX1 U34 ( .A(n1740), .B(n2036), .C(n600), .Z(n1741) );
  IVSVTX0H U35 ( .A(n356), .Z(n1780) );
  IVSVTX0H U36 ( .A(n1614), .Z(n1432) );
  IVSVTX2 U37 ( .A(n2077), .Z(n1678) );
  IVSVTX0H U38 ( .A(n570), .Z(n1431) );
  AO7SVTX1 U39 ( .A(n1501), .B(n1636), .C(n1461), .Z(n1502) );
  AO7SVTX1 U40 ( .A(n1694), .B(n1954), .C(n653), .Z(n1955) );
  ND2SVTX6 U41 ( .A(n1913), .B(n1920), .Z(n641) );
  EOSVTX0H U42 ( .A(n1449), .B(n1448), .Z(n789) );
  CTIVSVTX2 U43 ( .A(n260), .Z(n343) );
  NR2ASVTX1 U44 ( .A(n171), .B(n44), .Z(n603) );
  IVSVTX4 U45 ( .A(n175), .Z(n560) );
  IVSVTX0H U46 ( .A(n245), .Z(n1578) );
  AO7SVTX1 U47 ( .A(n182), .B(n1453), .C(n1589), .Z(n1590) );
  BFSVTX0H U48 ( .A(n1756), .Z(n1757) );
  IVSVTX0H U49 ( .A(n1870), .Z(n1778) );
  IVSVTX0H U50 ( .A(n1839), .Z(n110) );
  IVSVTX0H U51 ( .A(n1857), .Z(n1858) );
  IVSVTX0H U52 ( .A(n2049), .Z(n2050) );
  IVSVTX0H U53 ( .A(n2056), .Z(n2023) );
  IVSVTX0H U54 ( .A(n1944), .Z(n2058) );
  IVSVTX0H U55 ( .A(n1754), .Z(n1755) );
  IVSVTX0H U56 ( .A(n1840), .Z(n1841) );
  IVSVTX0H U57 ( .A(n1951), .Z(n1953) );
  IVSVTX0H U58 ( .A(n1881), .Z(n693) );
  IVSVTX0H U59 ( .A(n2015), .Z(n2016) );
  BFSVTX2 U60 ( .A(n1675), .Z(n2080) );
  IVSVTX0H U61 ( .A(n595), .Z(n1793) );
  IVSVTX0H U62 ( .A(n1864), .Z(n1865) );
  IVSVTX0H U63 ( .A(n683), .Z(n762) );
  IVSVTX0H U64 ( .A(n1941), .Z(n2019) );
  IVSVTX0H U65 ( .A(n1928), .Z(n1998) );
  IVSVTX0H U66 ( .A(n217), .Z(n1776) );
  IVSVTX0H U67 ( .A(n2037), .Z(n2038) );
  IVSVTX0H U68 ( .A(n1580), .Z(n1437) );
  NR2ASVTX1 U69 ( .A(n1958), .B(n1957), .Z(n1963) );
  IVSVTX0H U70 ( .A(n2017), .Z(n2018) );
  CTBUFSVTX8 U71 ( .A(n1575), .Z(n260) );
  IVSVTX0H U72 ( .A(n1969), .Z(n1705) );
  BFSVTX2 U73 ( .A(n43), .Z(n174) );
  IVSVTX0H U74 ( .A(n182), .Z(n1591) );
  ENSVTX0H U75 ( .A(n1752), .B(n231), .Z(n1753) );
  ND3SVTX4 U76 ( .A(n136), .B(n993), .C(n992), .Z(n1538) );
  B_ND2SVTX0H U77 ( .A(n1663), .B(n588), .Z(n1666) );
  NR2ASVTX1 U78 ( .A(n1124), .B(n44), .Z(n601) );
  IVSVTX0H U79 ( .A(n3), .Z(n1869) );
  NR2ASVTX2 U80 ( .A(m1[8]), .B(n44), .Z(n598) );
  ND2ASVTX4 U81 ( .A(n1390), .B(n1389), .Z(n1856) );
  IVSVTX2 U82 ( .A(n1375), .Z(n2040) );
  ND2SVTX8 U83 ( .A(n193), .B(n82), .Z(n406) );
  IVSVTX0H U84 ( .A(n1490), .Z(n1491) );
  IVSVTX0H U85 ( .A(n1727), .Z(n1498) );
  IVSVTX0H U86 ( .A(n1376), .Z(n1377) );
  IVSVTX0H U87 ( .A(n1885), .Z(n1984) );
  IVSVTX0H U88 ( .A(n1440), .Z(n1442) );
  IVSVTX0H U89 ( .A(n1374), .Z(n1375) );
  IVSVTX0H U90 ( .A(n1579), .Z(n1582) );
  IVSVTX0H U91 ( .A(n1814), .Z(n1815) );
  IVSVTX0H U92 ( .A(n1372), .Z(n1373) );
  ND2SVTX2 U93 ( .A(n57), .B(n1550), .Z(n668) );
  IVSVTX0H U94 ( .A(n1983), .Z(n1887) );
  IVSVTX0H U95 ( .A(n1884), .Z(n1986) );
  IVSVTX0H U96 ( .A(n190), .Z(n1829) );
  IVSVTX2 U97 ( .A(n1873), .Z(n1636) );
  CTIVSVTX2 U98 ( .A(n1567), .Z(n613) );
  IVSVTX0H U99 ( .A(n1300), .Z(n1147) );
  NR2ASVTX1 U100 ( .A(n218), .B(n297), .Z(n298) );
  IVSVTX0H U101 ( .A(n1927), .Z(n658) );
  IVSVTX0H U102 ( .A(n1758), .Z(n1760) );
  IVSVTX0H U103 ( .A(n1501), .Z(n1603) );
  ND2SVTX4 U104 ( .A(n583), .B(n1245), .Z(n1896) );
  IVSVTX0H U105 ( .A(n1782), .Z(n1872) );
  ND3ASVTX6 U106 ( .A(n316), .B(n315), .C(n313), .Z(n312) );
  IVSVTX0H U107 ( .A(n1759), .Z(n545) );
  IVSVTX4 U108 ( .A(n1165), .Z(n1568) );
  IVSVTX0H U109 ( .A(n1334), .Z(n1750) );
  AO7SVTX1 U110 ( .A(n672), .B(n1033), .C(n989), .Z(n990) );
  IVSVTX2 U111 ( .A(n757), .Z(n57) );
  IVSVTX0H U112 ( .A(n1820), .Z(n1737) );
  ND3SVTX4 U113 ( .A(n1421), .B(n1422), .C(n1420), .Z(n359) );
  NR2SVTX2 U114 ( .A(n1494), .B(n1493), .Z(n1727) );
  ND2ASVTX6 U115 ( .A(n938), .B(n167), .Z(n1429) );
  NR2ASVTX1 U116 ( .A(n515), .B(m1[24]), .Z(n989) );
  IVSVTX2 U117 ( .A(n1396), .Z(n2046) );
  IVSVTX0H U118 ( .A(n1735), .Z(n1819) );
  BFSVTX0H U119 ( .A(n1128), .Z(n138) );
  NR2SVTX4 U120 ( .A(n1243), .B(n1244), .Z(n1245) );
  ND2SVTX2 U121 ( .A(n822), .B(n1297), .Z(n997) );
  AO21DSVTX4 U122 ( .A(n1150), .B(n59), .C(n1416), .D(n1300), .Z(n1153) );
  AO6SVTX6 U123 ( .A(n58), .B(n729), .C(n1149), .Z(n1152) );
  AO7SVTX4 U124 ( .A(n722), .B(n719), .C(n1364), .Z(n1672) );
  AO7SVTX4 U125 ( .A(n436), .B(n266), .C(n1912), .Z(n265) );
  ND2SVTX2 U126 ( .A(n150), .B(n1482), .Z(n572) );
  IVSVTX8 U127 ( .A(n949), .Z(n1461) );
  IVSVTX2 U128 ( .A(n1150), .Z(n729) );
  IVSVTX2 U129 ( .A(n483), .Z(n757) );
  ND2ASVTX4 U130 ( .A(n1164), .B(n1277), .Z(n1912) );
  IVSVTX4 U131 ( .A(n1163), .Z(n266) );
  ND4ABSVTX6 U132 ( .A(n1241), .B(n9), .C(n1214), .D(n1213), .Z(n1210) );
  IVSVTX2 U133 ( .A(n34), .Z(n37) );
  AO4SVTX4 U134 ( .A(n194), .B(n1907), .C(n475), .D(n476), .Z(n470) );
  F_ND2ASVTX2 U135 ( .A(n1330), .B(n42), .Z(n1569) );
  NR2SVTX2 U136 ( .A(n1330), .B(n503), .Z(n483) );
  IVSVTX2 U137 ( .A(n60), .Z(n585) );
  ND3ASVTX4 U138 ( .A(n1296), .B(n1877), .C(n1303), .Z(n295) );
  IVSVTX6 U139 ( .A(n335), .Z(n195) );
  ND2ASVTX6 U140 ( .A(n34), .B(n478), .Z(n474) );
  IVSVTX0H U141 ( .A(n878), .Z(n820) );
  IVSVTX0H U142 ( .A(n1282), .Z(n1283) );
  ND2SVTX2 U143 ( .A(n503), .B(n488), .Z(n487) );
  F_ND2ASVTX2 U144 ( .A(n1323), .B(n1276), .Z(n1164) );
  AO21SVTX4 U145 ( .A(n240), .B(n1011), .C(n353), .D(n1016), .Z(n998) );
  ND2SVTX2 U146 ( .A(n472), .B(n1904), .Z(n476) );
  NR2SVTX2 U147 ( .A(n311), .B(n710), .Z(n202) );
  IVSVTX4 U148 ( .A(n60), .Z(n2036) );
  NR2SVTX2 U149 ( .A(n363), .B(n206), .Z(n205) );
  F_ND2ASVTX2 U150 ( .A(n210), .B(n1640), .Z(n1361) );
  OR3SVTX4 U151 ( .A(n1226), .B(n1220), .C(n1877), .Z(n802) );
  IVSVTX6 U152 ( .A(n34), .Z(n36) );
  CTIVSVTX6 U153 ( .A(n1601), .Z(n599) );
  BFSVTX10 U154 ( .A(n503), .Z(n591) );
  IVSVTX6 U155 ( .A(n41), .Z(n335) );
  BFSVTX4 U156 ( .A(n1558), .Z(n1559) );
  IVSVTX2 U157 ( .A(n963), .Z(n643) );
  IVSVTX0H U158 ( .A(n1286), .Z(n1287) );
  BFSVTX8 U159 ( .A(n1302), .Z(n1276) );
  CTIVSVTX2 U160 ( .A(n1556), .Z(n573) );
  ND2ASVTX4 U161 ( .A(n1978), .B(n1198), .Z(n1200) );
  ND2SVTX2 U162 ( .A(n1758), .B(n1360), .Z(n392) );
  NR2ASVTX2 U163 ( .A(n1903), .B(n1902), .Z(n1905) );
  F_ENSVTX2 U164 ( .A(n1208), .B(n40), .Z(n464) );
  CTIVSVTX2 U165 ( .A(n753), .Z(n1342) );
  IVSVTX0H U166 ( .A(n1177), .Z(n362) );
  BFSVTX4 U167 ( .A(n1009), .Z(n1033) );
  IVSVTX0H U168 ( .A(n1255), .Z(n1260) );
  IVSVTX2 U169 ( .A(n735), .Z(n706) );
  BFSVTX8 U170 ( .A(n811), .Z(n495) );
  ND2ASVTX6 U171 ( .A(n59), .B(n1553), .Z(n1031) );
  IVSVTX0H U172 ( .A(n1067), .Z(n308) );
  IVSVTX0H U173 ( .A(n1331), .Z(n1333) );
  NR2SVTX2 U174 ( .A(n1063), .B(n311), .Z(n262) );
  F_ND2ASVTX2 U175 ( .A(n73), .B(n1359), .Z(n1360) );
  IVSVTX4 U176 ( .A(n578), .Z(n1251) );
  IVSVTX4 U177 ( .A(n43), .Z(n1902) );
  NR2ASVTX2 U178 ( .A(n961), .B(n390), .Z(n645) );
  AO2SVTX6 U179 ( .A(n449), .B(n448), .C(n1756), .D(n1330), .Z(n447) );
  BFSVTX6 U180 ( .A(n1978), .Z(n60) );
  ND4SVTX6 U181 ( .A(n1640), .B(n1059), .C(n1057), .D(n1058), .Z(n334) );
  NR2SVTX2 U182 ( .A(n1075), .B(n746), .Z(n497) );
  NR2ASVTX1 U183 ( .A(n1172), .B(n1171), .Z(n1176) );
  ND2SVTX1 U184 ( .A(n1177), .B(n1171), .Z(n1170) );
  ND2ASVTX4 U185 ( .A(n1038), .B(n1043), .Z(n714) );
  IVSVTX6 U186 ( .A(n1337), .Z(n1339) );
  IVSVTX6 U187 ( .A(n231), .Z(n232) );
  CTIVSVTX4 U188 ( .A(n317), .Z(n514) );
  IVSVTX6 U189 ( .A(n38), .Z(n39) );
  ND2SVTX2 U190 ( .A(n364), .B(n371), .Z(n756) );
  IVSVTX0H U191 ( .A(n916), .Z(n1203) );
  ND2ASVTX6 U192 ( .A(n425), .B(n424), .Z(n1014) );
  CTIVSVTX2 U193 ( .A(n451), .Z(n146) );
  IVSVTX8 U194 ( .A(n1248), .Z(n1435) );
  IVSVTX2 U195 ( .A(n1072), .Z(n499) );
  NR2SVTX2 U196 ( .A(n1065), .B(n1062), .Z(n1063) );
  NR3SVTX6 U197 ( .A(n649), .B(n1160), .C(n1159), .Z(n648) );
  ND2SVTX6 U198 ( .A(n1310), .B(n317), .Z(n1543) );
  IVSVTX2 U199 ( .A(n1011), .Z(n1012) );
  IVSVTX0H U200 ( .A(n1173), .Z(n1174) );
  AO6ABSVTX4 U201 ( .A(n981), .B(n1181), .C(n982), .Z(n983) );
  ND3SVTX6 U202 ( .A(n1039), .B(n1042), .C(n710), .Z(n1045) );
  IVSVTX4 U203 ( .A(n34), .Z(n35) );
  ND2SVTX2 U204 ( .A(n968), .B(n967), .Z(n247) );
  AO3NSVTX4 U205 ( .A(n231), .B(n1028), .C(n1026), .D(n1027), .Z(n795) );
  AO7NSVTX4 U206 ( .A(n1156), .B(n1158), .C(n872), .Z(n801) );
  NR2ASVTX2 U207 ( .A(n178), .B(n1034), .Z(n991) );
  ND2SVTX8 U208 ( .A(n1046), .B(n63), .Z(n1171) );
  IVSVTX6 U209 ( .A(n1320), .Z(n1248) );
  IVSVTX2 U210 ( .A(n517), .Z(n581) );
  IVSVTX2 U211 ( .A(n1080), .Z(n433) );
  IVSVTX0H U212 ( .A(n1079), .Z(n1024) );
  NR2SVTX2 U213 ( .A(n1042), .B(n1043), .Z(n125) );
  F_AN2SVTX2 U214 ( .A(n1000), .B(n78), .Z(n999) );
  NR2SVTX2 U215 ( .A(n47), .B(n46), .Z(n119) );
  IVSVTX2 U216 ( .A(n569), .Z(n568) );
  ND2SVTX2 U217 ( .A(n1169), .B(n1173), .Z(n960) );
  IVSVTX2 U218 ( .A(n818), .Z(n967) );
  IVSVTX0H U219 ( .A(n965), .Z(n966) );
  BFSVTX4 U220 ( .A(n1181), .Z(n166) );
  IVSVTX2 U221 ( .A(n1355), .Z(n67) );
  IVSVTX6 U222 ( .A(n519), .Z(n539) );
  IVSVTX2 U223 ( .A(n961), .Z(n46) );
  IVSVTX0H U224 ( .A(n981), .Z(n1180) );
  IVSVTX4 U225 ( .A(n1040), .Z(n1043) );
  IVSVTX2 U226 ( .A(n887), .Z(n1065) );
  AO7SVTX1 U227 ( .A(n965), .B(n506), .C(n964), .Z(n969) );
  ND2SVTX4 U228 ( .A(n818), .B(n427), .Z(n366) );
  BFSVTX2 U229 ( .A(n556), .Z(n127) );
  ND2SVTX2 U230 ( .A(n1414), .B(n1189), .Z(n574) );
  IVSVTX10 U231 ( .A(n479), .Z(n43) );
  IVSVTX0H U232 ( .A(n1169), .Z(n651) );
  IVSVTX6 U233 ( .A(n178), .Z(n672) );
  ND2ASVTX4 U234 ( .A(n72), .B(n252), .Z(n251) );
  IVSVTX8 U235 ( .A(n233), .Z(n231) );
  BFSVTX4 U236 ( .A(n83), .Z(n178) );
  ND2ASVTX6 U237 ( .A(n927), .B(n926), .Z(n491) );
  B_ND2SVTX2 U238 ( .A(n1142), .B(n296), .Z(n1312) );
  IVSVTX2 U239 ( .A(n707), .Z(n853) );
  ND2SVTX4 U240 ( .A(n517), .B(n911), .Z(n914) );
  CTIVSVTX2 U241 ( .A(n680), .Z(n774) );
  B_ND2SVTX2 U242 ( .A(n995), .B(n994), .Z(n961) );
  ND2SVTX6 U243 ( .A(n1587), .B(n1313), .Z(n1623) );
  ND2ASVTX4 U244 ( .A(n1306), .B(n1659), .Z(n252) );
  IVSVTX2 U245 ( .A(n1145), .Z(n1308) );
  F_ND2ASVTX2 U246 ( .A(n75), .B(n854), .Z(n372) );
  NR2SVTX1 U247 ( .A(m1[23]), .B(n1082), .Z(n23) );
  EN3SVTX6 U248 ( .A(n1126), .B(n347), .C(n79), .Z(n1090) );
  IVSVTX2 U249 ( .A(n1179), .Z(n982) );
  NR2ASVTX6 U250 ( .A(n775), .B(n65), .Z(n426) );
  ND2SVTX4 U251 ( .A(n1060), .B(n887), .Z(n680) );
  IVSVTX2 U252 ( .A(n542), .Z(n520) );
  IVSVTX2 U253 ( .A(n588), .Z(n685) );
  NR2ASVTX2 U254 ( .A(n928), .B(m1[24]), .Z(n1086) );
  IVSVTX2 U255 ( .A(n1305), .Z(n1306) );
  ND2SVTX2 U256 ( .A(n632), .B(n1271), .Z(n870) );
  CTIVSVTX4 U257 ( .A(n920), .Z(n320) );
  ND2SVTX4 U258 ( .A(n294), .B(n400), .Z(n1305) );
  ND2SVTX2 U259 ( .A(n953), .B(n294), .Z(n1247) );
  AN2SVTX2 U260 ( .A(n481), .B(m1[23]), .Z(n788) );
  NR2SVTX4 U261 ( .A(n1450), .B(n747), .Z(n213) );
  IVSVTX2 U262 ( .A(n666), .Z(n96) );
  ND2ASVTX6 U263 ( .A(n85), .B(n79), .Z(n1346) );
  ND2ASVTX6 U264 ( .A(n423), .B(n354), .Z(n1758) );
  ND2SVTX2 U265 ( .A(n99), .B(m1[20]), .Z(n1184) );
  BFSVTX6 U266 ( .A(n1664), .Z(n508) );
  ND2ASVTX4 U267 ( .A(n953), .B(n83), .Z(n1179) );
  ND2SVTX2 U268 ( .A(n708), .B(n154), .Z(n1318) );
  IVSVTX6 U269 ( .A(n1659), .Z(n64) );
  NR2SVTX6 U270 ( .A(n851), .B(n1299), .Z(n919) );
  ND2SVTX4 U271 ( .A(n1820), .B(n740), .Z(n1501) );
  NR2SVTX6 U272 ( .A(n949), .B(n403), .Z(n402) );
  NR3SVTX6 U273 ( .A(m1[23]), .B(n211), .C(n294), .Z(n775) );
  IVSVTX4 U274 ( .A(n964), .Z(n1299) );
  ND2ASVTX6 U275 ( .A(m1[20]), .B(n1068), .Z(n886) );
  IVSVTX6 U276 ( .A(n83), .Z(n556) );
  IVSVTX2 U277 ( .A(n1632), .Z(n749) );
  NR2ASVTX4 U278 ( .A(m1[14]), .B(m1[16]), .Z(n245) );
  NR2SVTX4 U279 ( .A(n928), .B(m1[24]), .Z(n980) );
  CTIVSVTX2 U280 ( .A(n85), .Z(n709) );
  CTIVSVTX2 U281 ( .A(n616), .Z(n852) );
  IVSVTX2 U282 ( .A(n84), .Z(n444) );
  ND2SVTX4 U283 ( .A(n842), .B(n841), .Z(n1257) );
  ND2SVTX4 U284 ( .A(n1494), .B(n1493), .Z(n292) );
  IVSVTX2 U285 ( .A(n1288), .Z(n826) );
  NR2SVTX6 U286 ( .A(n1580), .B(n509), .Z(n1664) );
  AN2SVTX4 U287 ( .A(n1000), .B(n964), .Z(n239) );
  ND2SVTX6 U288 ( .A(n695), .B(n696), .Z(n1681) );
  NR2SVTX2 U289 ( .A(n1734), .B(n1733), .Z(n740) );
  ND2SVTX4 U290 ( .A(n1663), .B(n1317), .Z(n1355) );
  IVSVTX6 U291 ( .A(n75), .Z(n605) );
  ND2ASVTX6 U292 ( .A(m1[16]), .B(n347), .Z(n712) );
  ND2ASVTX4 U293 ( .A(n752), .B(n400), .Z(n952) );
  IVSVTX2 U294 ( .A(n619), .Z(n1137) );
  ND2ASVTX6 U295 ( .A(n410), .B(n82), .Z(n1474) );
  IVSVTX2 U296 ( .A(n1096), .Z(n695) );
  IVSVTX6 U297 ( .A(n760), .Z(n761) );
  NR3SVTX4 U298 ( .A(n816), .B(n347), .C(n617), .Z(n844) );
  IVSVTX8 U299 ( .A(n1068), .Z(n76) );
  IVSVTX4 U300 ( .A(n167), .Z(n154) );
  NR2SVTX4 U301 ( .A(n586), .B(n1399), .Z(n428) );
  IVSVTX2 U302 ( .A(n1138), .Z(n71) );
  IVSVTX4 U303 ( .A(n1194), .Z(n49) );
  ND2ASVTX4 U304 ( .A(m1[17]), .B(n400), .Z(n399) );
  IVSVTX2 U305 ( .A(n1384), .Z(n1111) );
  ND2ASVTX4 U306 ( .A(m1[20]), .B(n75), .Z(n1169) );
  ND2SVTX6 U307 ( .A(n1125), .B(n543), .Z(n1494) );
  F_ND2ASVTX2 U308 ( .A(n1123), .B(n504), .Z(n1100) );
  IVSVTX6 U309 ( .A(n752), .Z(n89) );
  ND2ASVTX4 U310 ( .A(m1[8]), .B(n259), .Z(n1862) );
  IVSVTX8 U311 ( .A(n346), .Z(n347) );
  ND2ASVTX6 U312 ( .A(n752), .B(n193), .Z(n1428) );
  F_IVSVTX1 U313 ( .A(n708), .Z(n86) );
  IVSVTX10 U314 ( .A(n743), .Z(n1068) );
  CTIVSVTX6 U315 ( .A(n226), .Z(n79) );
  IVSVTX6 U316 ( .A(n928), .Z(n507) );
  IVSVTX2 U317 ( .A(n857), .Z(n140) );
  IVSVTX2 U318 ( .A(n1733), .Z(n258) );
  ND2SVTX2 U319 ( .A(m1[8]), .B(n1106), .Z(n1959) );
  B_ND2SVTX2 U320 ( .A(n1093), .B(n1092), .Z(n1384) );
  IVSVTX4 U321 ( .A(n52), .Z(n528) );
  ND2ASVTX4 U322 ( .A(n752), .B(n171), .Z(n1579) );
  AO7SVTX4 U323 ( .A(n1116), .B(n299), .C(n738), .Z(n1104) );
  AO7SVTX6 U324 ( .A(n653), .B(n1951), .C(n1952), .Z(n1864) );
  NR2SVTX6 U325 ( .A(n84), .B(n1479), .Z(n566) );
  NR2SVTX4 U326 ( .A(n1995), .B(n1928), .Z(n942) );
  AO6ABSVTX4 U327 ( .A(n1786), .B(n765), .C(n907), .Z(n908) );
  ND2SVTX2 U328 ( .A(n816), .B(n1519), .Z(n1996) );
  AO7SVTX4 U329 ( .A(m1[16]), .B(n889), .C(n752), .Z(n224) );
  CTIVSVTX6 U330 ( .A(n410), .Z(n526) );
  IVSVTX8 U331 ( .A(n1345), .Z(n48) );
  IVSVTX2 U332 ( .A(n950), .Z(n87) );
  CTIVSVTX4 U333 ( .A(n617), .Z(n463) );
  NR2SVTX6 U334 ( .A(n759), .B(n752), .Z(n1733) );
  IVSVTX2 U335 ( .A(n728), .Z(n357) );
  IVSVTX8 U336 ( .A(n743), .Z(n744) );
  IVSVTX2 U337 ( .A(n835), .Z(n2044) );
  ND2SVTX2 U338 ( .A(n259), .B(n752), .Z(n546) );
  NR2SVTX6 U339 ( .A(m1[12]), .B(n462), .Z(n1734) );
  ND2ASVTX4 U340 ( .A(n906), .B(n938), .Z(n1801) );
  NR2SVTX4 U341 ( .A(n1519), .B(n896), .Z(n2024) );
  ND2SVTX2 U342 ( .A(m1[16]), .B(n889), .Z(n225) );
  IVSVTX4 U343 ( .A(n861), .Z(n1370) );
  ND2SVTX6 U344 ( .A(n90), .B(n654), .Z(n653) );
  NR2SVTX4 U345 ( .A(n1792), .B(n1102), .Z(n1957) );
  IVSVTX6 U346 ( .A(m1[27]), .Z(n608) );
  IVSVTX4 U347 ( .A(n430), .Z(n192) );
  AO7SVTX4 U348 ( .A(n1983), .B(n1881), .C(n1882), .Z(n904) );
  IVSVTX6 U349 ( .A(n906), .Z(n1124) );
  ND2ASVTX4 U350 ( .A(m1[10]), .B(m1[12]), .Z(n1828) );
  ND2ASVTX4 U351 ( .A(n1792), .B(n713), .Z(n728) );
  ND2SVTX4 U352 ( .A(n1123), .B(n758), .Z(n950) );
  CTIVSVTX4 U353 ( .A(n2003), .Z(n80) );
  IVSVTX6 U354 ( .A(n944), .Z(n1102) );
  IVSVTX6 U355 ( .A(n860), .Z(n307) );
  ND2ASVTX6 U356 ( .A(n155), .B(n895), .Z(n1524) );
  ND2SVTX4 U357 ( .A(m1[8]), .B(n898), .Z(n861) );
  IVSVTX10 U358 ( .A(n1126), .Z(n1345) );
  OR2BSVTX6 U359 ( .A(m1[1]), .B(m1[4]), .Z(n1529) );
  ND2ASVTX6 U360 ( .A(n906), .B(n713), .Z(n1827) );
  ND3ASVTX6 U361 ( .A(m1[0]), .B(n758), .C(n939), .Z(n617) );
  CTBUFSVTX8 U362 ( .A(m1[2]), .Z(n1934) );
  NR2SVTX2 U363 ( .A(m1[10]), .B(n751), .Z(n1723) );
  IVSVTX6 U364 ( .A(n743), .Z(n760) );
  NR2ASVTX4 U365 ( .A(n733), .B(m1[12]), .Z(n386) );
  IVSVTX2 U366 ( .A(n1367), .Z(n10) );
  ND2SVTX6 U367 ( .A(n243), .B(m1[17]), .Z(n1612) );
  IVSVTX4 U368 ( .A(n675), .Z(n446) );
  IVSVTX6 U369 ( .A(m1[23]), .Z(n93) );
  NR3SVTX4 U370 ( .A(n896), .B(n160), .C(n2004), .Z(n268) );
  IVSVTX8 U371 ( .A(n1792), .Z(n654) );
  AO7SVTX2 U372 ( .A(n91), .B(n297), .C(n939), .Z(n271) );
  ND2ASVTX4 U373 ( .A(m1[17]), .B(n430), .Z(n1647) );
  NR3ABSVTX4 U374 ( .A(n1123), .B(n898), .C(n20), .Z(n208) );
  IVSVTX10 U375 ( .A(m1[17]), .Z(n1126) );
  IVSVTX10 U376 ( .A(n951), .Z(n889) );
  IVSVTX10 U377 ( .A(n751), .Z(n938) );
  BFSVTX8 U378 ( .A(n733), .Z(n297) );
  IVSVTX6 U379 ( .A(n1130), .Z(n855) );
  IVSVTX10 U380 ( .A(n346), .Z(n1131) );
  IVSVTX10 U381 ( .A(n244), .Z(n82) );
  IVSVTX8 U382 ( .A(n1106), .Z(n122) );
  IVSVTX8 U383 ( .A(n894), .Z(n738) );
  IVSVTX4 U384 ( .A(n1094), .Z(n1975) );
  ND3SVTX4 U385 ( .A(n218), .B(m1[1]), .C(n734), .Z(n272) );
  F_ND2ASVTX2 U386 ( .A(n273), .B(n299), .Z(n2003) );
  IVSVTX10 U387 ( .A(n750), .Z(n751) );
  IVSVTX10 U388 ( .A(m1[8]), .Z(n860) );
  BFSVTX12 U389 ( .A(m1[0]), .Z(n218) );
  IVSVTX6 U390 ( .A(n733), .Z(n299) );
  IVSVTX6 U391 ( .A(m1[10]), .Z(n482) );
  IVSVTX4 U392 ( .A(m1[6]), .Z(n273) );
  NR2SVTX2 U393 ( .A(n1519), .B(m1[1]), .Z(n1932) );
  NR2ASVTX4 U394 ( .A(n472), .B(n1908), .Z(n194) );
  AO7SVTX2 U395 ( .A(n1105), .B(n1775), .C(n1124), .Z(n1098) );
  ND3SVTX4 U396 ( .A(n1914), .B(n640), .C(n641), .Z(n639) );
  NR2SVTX2 U397 ( .A(n515), .B(n1601), .Z(n848) );
  B_ND2SVTX2 U398 ( .A(n1344), .B(n1345), .Z(n1362) );
  IVSVTX8 U399 ( .A(n1207), .Z(n38) );
  IVSVTX10 U400 ( .A(m1[2]), .Z(n896) );
  AO2SVTX6 U401 ( .A(n1019), .B(n1670), .C(n1018), .D(n1017), .Z(n454) );
  ND3ABSVTX6 U402 ( .A(n49), .B(n1261), .C(n355), .Z(n622) );
  IVSVTX4 U403 ( .A(n1141), .Z(n541) );
  ND2SVTX2 U404 ( .A(n279), .B(n471), .Z(n473) );
  ND2SVTX2 U405 ( .A(n1938), .B(n1385), .Z(n1386) );
  AO7SVTX4 U406 ( .A(n1625), .B(n1453), .C(n1624), .Z(n1626) );
  ND4SVTX8 U407 ( .A(n1510), .B(n1511), .C(n120), .D(n1513), .Z(m2[11]) );
  IVSVTX4 U408 ( .A(n121), .Z(n120) );
  AO2SVTX2 U409 ( .A(n2071), .B(n2070), .C(n174), .D(n2069), .Z(n2072) );
  ND2SVTX2 U410 ( .A(n174), .B(n1456), .Z(n1469) );
  F_ENSVTX2 U411 ( .A(n1607), .B(n1606), .Z(n1608) );
  F_EOSVTX2 U412 ( .A(n1619), .B(n1618), .Z(n1620) );
  AO6SVTX4 U413 ( .A(n219), .B(n1617), .C(n1616), .Z(n1618) );
  AO21SVTX4 U414 ( .A(n1636), .B(n1635), .C(n1501), .D(n1634), .Z(n1637) );
  AO7ABSVTX4 U415 ( .A(m1[10]), .B(m1[8]), .C(n505), .Z(n773) );
  IVSVTX4 U416 ( .A(n1452), .Z(n1453) );
  AO6SVTX6 U417 ( .A(n1885), .B(n905), .C(n904), .Z(n1788) );
  F_ENSVTX2 U418 ( .A(n1739), .B(n1738), .Z(n1740) );
  AO8SVTX2 U419 ( .A(n1597), .B(n1505), .C(n1870), .D(n1447), .Z(n1448) );
  ND2SVTX2 U420 ( .A(n14), .B(n66), .Z(n1635) );
  IVSVTX2 U421 ( .A(n187), .Z(n1625) );
  AO7ASVTX8 U422 ( .A(n43), .B(n1425), .C(n1424), .Z(n286) );
  ND2SVTX4 U423 ( .A(n1677), .B(n1676), .Z(n2076) );
  ENSVTX8 U424 ( .A(n1901), .B(n1900), .Z(m2[18]) );
  AO6CSVTX4 U425 ( .A(n233), .B(n1334), .C(n1751), .Z(n1335) );
  NR2SVTX4 U426 ( .A(n721), .B(n532), .Z(n628) );
  IVSVTX6 U427 ( .A(n318), .Z(n1336) );
  AO6SVTX8 U428 ( .A(n1646), .B(n827), .C(n1), .Z(n13) );
  AO7SVTX8 U429 ( .A(n1644), .B(n831), .C(n1641), .Z(n1) );
  IVSVTX8 U430 ( .A(n715), .Z(n716) );
  ENSVTX4 U431 ( .A(n814), .B(n1335), .Z(n554) );
  IVSVTX8 U432 ( .A(n715), .Z(n1519) );
  ND2SVTX8 U433 ( .A(n903), .B(n1368), .Z(n910) );
  IVSVTX8 U434 ( .A(n1115), .Z(n2062) );
  IVSVTX10 U435 ( .A(m1[3]), .Z(n733) );
  ND3ABSVTX6 U436 ( .A(n1902), .B(n672), .C(n1148), .Z(n1149) );
  AO7SVTX6 U437 ( .A(n1250), .B(n581), .C(n579), .Z(n578) );
  AO3SVTX8 U438 ( .A(n341), .B(n612), .C(n338), .D(n337), .Z(m2[25]) );
  BFSVTX1 U439 ( .A(n1777), .Z(n3) );
  AO7ABSVTX8 U440 ( .A(n1298), .B(n370), .C(n5), .Z(n1302) );
  AO7ABSVTX6 U441 ( .A(n840), .B(n883), .C(n642), .Z(n5) );
  ND3ASVTX8 U442 ( .A(m1[20]), .B(n852), .C(n157), .Z(n850) );
  ENSVTX8 U443 ( .A(n1000), .B(n533), .Z(n1019) );
  EO3SVTX8 U444 ( .A(n898), .B(n1106), .C(n734), .Z(n1113) );
  AO7SVTX4 U445 ( .A(n1056), .B(n1055), .C(n1054), .Z(n1057) );
  AO1ASVTX8 U446 ( .A(n6), .B(n662), .C(n660), .D(n659), .Z(m2[22]) );
  IVSVTX4 U447 ( .A(n8), .Z(n1053) );
  ND2SVTX4 U448 ( .A(n1049), .B(n1173), .Z(n8) );
  IVSVTX4 U449 ( .A(n244), .Z(n430) );
  IVSVTX4 U450 ( .A(n739), .Z(n66) );
  AO1ASVTX6 U451 ( .A(n181), .B(n622), .C(n1200), .D(n621), .Z(n9) );
  IVSVTX10 U452 ( .A(n817), .Z(n1116) );
  AO6SVTX8 U453 ( .A(n1430), .B(n1351), .C(n1350), .Z(n489) );
  IVSVTX8 U454 ( .A(n944), .Z(n1105) );
  IVSVTX4 U455 ( .A(n51), .Z(n1687) );
  NR2ASVTX6 U456 ( .A(n51), .B(n10), .Z(n1884) );
  ND2SVTX4 U457 ( .A(n894), .B(m1[8]), .Z(n51) );
  AO7SVTX6 U458 ( .A(n909), .B(n1788), .C(n908), .Z(n717) );
  AO7SVTX6 U459 ( .A(n2039), .B(n1370), .C(n1371), .Z(n862) );
  ND2SVTX4 U460 ( .A(n1116), .B(n860), .Z(n1371) );
  IVSVTX4 U461 ( .A(n45), .Z(n42) );
  NR2ASVTX6 U462 ( .A(n45), .B(n554), .Z(n550) );
  IVSVTX8 U463 ( .A(n1357), .Z(n41) );
  ND2ASVTX8 U464 ( .A(n1109), .B(n1107), .Z(n1115) );
  IVSVTX10 U465 ( .A(m1[12]), .Z(n410) );
  ND2SVTX4 U466 ( .A(n452), .B(n43), .Z(n451) );
  NR4ABCSVTX8 U467 ( .A(n77), .B(n381), .C(n761), .D(n616), .Z(n460) );
  IVSVTX10 U468 ( .A(n167), .Z(n193) );
  ND2SVTX4 U469 ( .A(n1722), .B(n11), .Z(n830) );
  ND2SVTX4 U470 ( .A(n204), .B(n1721), .Z(n11) );
  ND2ASVTX8 U471 ( .A(n759), .B(n82), .Z(n1721) );
  ND2SVTX6 U472 ( .A(n421), .B(n420), .Z(n1319) );
  ND3SVTX8 U473 ( .A(n639), .B(n637), .C(n636), .Z(m2[20]) );
  ND2SVTX6 U474 ( .A(n19), .B(n558), .Z(n692) );
  BFSVTX4 U475 ( .A(n1674), .Z(n1677) );
  IVSVTX8 U476 ( .A(n951), .Z(n1130) );
  ND2ASVTX8 U477 ( .A(n1138), .B(n619), .Z(n1141) );
  IVSVTX4 U478 ( .A(n97), .Z(n114) );
  BFSVTX10 U479 ( .A(n752), .Z(n12) );
  ND3SVTX4 U480 ( .A(n398), .B(n524), .C(n401), .Z(n397) );
  AO7SVTX8 U481 ( .A(n300), .B(n1651), .C(n13), .Z(n230) );
  BFSVTX1 U482 ( .A(n1632), .Z(n14) );
  AO20SVTX8 U483 ( .A(n15), .B(n1008), .C(n36), .D(n1007), .Z(n1550) );
  IVSVTX4 U484 ( .A(n16), .Z(n15) );
  AO7SVTX6 U485 ( .A(n1006), .B(n1005), .C(n1000), .Z(n16) );
  MUX21NSVTX8 U486 ( .A(n392), .B(n1360), .S(n391), .Z(n544) );
  AO7SVTX8 U487 ( .A(n1840), .B(n1837), .C(n1838), .Z(n1495) );
  ND2ASVTX8 U488 ( .A(n291), .B(n1134), .Z(n1840) );
  EOSVTX8 U489 ( .A(n999), .B(n306), .Z(n1003) );
  BFSVTX1 U490 ( .A(n1647), .Z(n17) );
  AO6SVTX8 U491 ( .A(n1430), .B(n1307), .C(n251), .Z(n250) );
  IVSVTX12 U492 ( .A(n38), .Z(n40) );
  IVSVTX8 U493 ( .A(n884), .Z(n885) );
  ND2SVTX4 U494 ( .A(n482), .B(n856), .Z(n1952) );
  BFSVTX1 U495 ( .A(n1769), .Z(n18) );
  IVSVTX4 U496 ( .A(n393), .Z(n19) );
  IVSVTX4 U497 ( .A(n860), .Z(n20) );
  IVSVTX2 U498 ( .A(n1055), .Z(n1052) );
  ND2SVTX4 U499 ( .A(m1[24]), .B(n76), .Z(n1060) );
  IVSVTX2 U500 ( .A(n61), .Z(n358) );
  IVSVTX4 U501 ( .A(n1314), .Z(n289) );
  F_MUX21NSVTX1 U502 ( .A(n1256), .B(n1262), .S(n1255), .Z(n1258) );
  AN2SVTX0H U503 ( .A(n840), .B(n882), .Z(n783) );
  F_ND2SVTX0H U504 ( .A(n150), .B(n1479), .Z(n1484) );
  IVSVTX2 U505 ( .A(m1[24]), .Z(n240) );
  IVSVTX4 U506 ( .A(n1142), .Z(n748) );
  IVSVTX2 U507 ( .A(n731), .Z(n732) );
  BFSVTX1 U508 ( .A(n2011), .Z(n2065) );
  NR2ASVTX1 U509 ( .A(n259), .B(n44), .Z(n600) );
  AO17SVTX2 U510 ( .A(n1548), .B(n1549), .C(n1547), .D(n43), .Z(n437) );
  F_ND2SVTX0H U511 ( .A(n1681), .B(n1682), .Z(n1686) );
  F_ND2SVTX0H U512 ( .A(n1475), .B(n1474), .Z(n1478) );
  NR2ASVTX1 U513 ( .A(n1587), .B(n541), .Z(n1593) );
  NR2ASVTX1 U514 ( .A(n526), .B(n44), .Z(n602) );
  F_ND2SVTX0H U515 ( .A(n2071), .B(n1892), .Z(n1893) );
  F_ND2SVTX0H U516 ( .A(n1509), .B(n37), .Z(n1510) );
  AN2SVTX6 U517 ( .A(n1305), .B(n712), .Z(n21) );
  AN2SVTX0H U518 ( .A(n2071), .B(n1993), .Z(n22) );
  IVSVTX10 U519 ( .A(n273), .Z(n90) );
  IVSVTX12 U520 ( .A(n744), .Z(n75) );
  IVSVTX12 U521 ( .A(m1[25]), .Z(n515) );
  ND2SVTX2 U522 ( .A(n1068), .B(n1000), .Z(n1061) );
  IVSVTX2 U523 ( .A(n851), .Z(n70) );
  IVSVTX12 U524 ( .A(m1[24]), .Z(n1000) );
  IVSVTX10 U525 ( .A(n99), .Z(n83) );
  IVSVTX6 U526 ( .A(m1[23]), .Z(n99) );
  IVSVTX10 U527 ( .A(n482), .Z(n462) );
  AO7SVTX6 U528 ( .A(n2017), .B(n2015), .C(n414), .Z(n1376) );
  IVSVTX12 U529 ( .A(n896), .Z(n816) );
  AN2SVTX4 U530 ( .A(n947), .B(n782), .Z(n24) );
  IVSVTX8 U531 ( .A(m1[20]), .Z(n953) );
  IVSVTX12 U532 ( .A(m1[20]), .Z(n226) );
  IVSVTX4 U533 ( .A(m1[20]), .Z(n481) );
  IVSVTX12 U534 ( .A(m1[16]), .Z(n167) );
  AN3SVTX6 U535 ( .A(n463), .B(n381), .C(n77), .Z(n25) );
  IVSVTX8 U536 ( .A(m1[19]), .Z(n346) );
  AN2SVTX0H U537 ( .A(n632), .B(n1270), .Z(n26) );
  AO7NSVTX4 U538 ( .A(n1458), .B(n1462), .C(n1457), .Z(n27) );
  IVSVTX4 U539 ( .A(n1658), .Z(n72) );
  IVSVTX12 U540 ( .A(n855), .Z(n171) );
  AO7NSVTX4 U541 ( .A(n65), .B(n369), .C(n1299), .Z(n28) );
  IVSVTX6 U542 ( .A(n163), .Z(n1227) );
  AO6SVTX8 U543 ( .A(n241), .B(n239), .C(n842), .Z(n163) );
  IVSVTX10 U544 ( .A(n1877), .Z(n45) );
  AN3SVTX4 U545 ( .A(n1601), .B(n1276), .C(n1188), .Z(n29) );
  AN2SVTX4 U546 ( .A(n387), .B(n1346), .Z(n30) );
  AO7ABSVTX8 U547 ( .A(n1276), .B(n1275), .C(n1274), .Z(n742) );
  AN3SVTX6 U548 ( .A(n870), .B(n1270), .C(n389), .Z(n31) );
  AO7NSVTX4 U549 ( .A(n458), .B(n41), .C(n184), .Z(n32) );
  NR2SVTX2 U550 ( .A(n473), .B(n618), .Z(n1909) );
  F_ND2SVTX1 U551 ( .A(n1850), .B(n1849), .Z(n1852) );
  ND2SVTX2 U552 ( .A(n1849), .B(n1850), .Z(n200) );
  AO4SVTX6 U553 ( .A(n1850), .B(n1849), .C(n1854), .D(n1853), .Z(n1122) );
  AO7CSVTX4 U554 ( .A(n127), .B(n1009), .C(m1[24]), .Z(n875) );
  IVSVTX12 U555 ( .A(n45), .Z(n34) );
  IVSVTX8 U556 ( .A(n1558), .Z(n62) );
  ND4ABSVTX8 U557 ( .A(n1569), .B(n1567), .C(n312), .D(n1568), .Z(n592) );
  F_ND2ASVTX2 U558 ( .A(n49), .B(n1255), .Z(n536) );
  AO7SVTX8 U559 ( .A(n142), .B(n1097), .C(n1682), .Z(n1855) );
  IVSVTX12 U560 ( .A(m1[7]), .Z(n944) );
  IVSVTX8 U561 ( .A(n1146), .Z(n1544) );
  IVSVTX12 U562 ( .A(m1[4]), .Z(n715) );
  IVSVTX6 U563 ( .A(n1327), .Z(n1451) );
  ND3SVTX4 U564 ( .A(n576), .B(n577), .C(n587), .Z(n302) );
  ND3SVTX4 U565 ( .A(n279), .B(n471), .C(n474), .Z(n468) );
  ND4SVTX6 U566 ( .A(n1950), .B(n1949), .C(n1948), .D(n1947), .Z(m2[1]) );
  AO2ABSVTX4 U567 ( .C(n2071), .D(n1846), .A(n1902), .B(n1845), .Z(n1847) );
  ND2SVTX6 U568 ( .A(n591), .B(n464), .Z(n1213) );
  F_ENSVTX2 U569 ( .A(n797), .B(n647), .Z(n1571) );
  F_ND2ASVTX2 U570 ( .A(n988), .B(n599), .Z(n993) );
  CTIVSVTX2 U571 ( .A(n1905), .Z(n475) );
  ND3SVTX4 U572 ( .A(n1237), .B(n573), .C(n706), .Z(n1212) );
  IVSVTX2 U573 ( .A(n754), .Z(n1023) );
  AO17SVTX4 U574 ( .A(n238), .B(n237), .C(n1288), .D(n1287), .Z(n1289) );
  AO7ASVTX6 U575 ( .A(n1203), .B(n1066), .C(n221), .Z(n918) );
  AO17SVTX4 U576 ( .A(n238), .B(n237), .C(n358), .D(n166), .Z(n1182) );
  AO7SVTX4 U577 ( .A(n1080), .B(n231), .C(n23), .Z(n754) );
  F_EOSVTX2 U578 ( .A(n1666), .B(n1665), .Z(n1667) );
  ND2ASVTX4 U579 ( .A(n1174), .B(n390), .Z(n1175) );
  F_ND2ASVTX2 U580 ( .A(n127), .B(n1542), .Z(n1546) );
  IVSVTX2 U581 ( .A(n793), .Z(n310) );
  AO7SVTX2 U582 ( .A(n1985), .B(n1834), .C(n1833), .Z(n1835) );
  CTIVSVTX2 U583 ( .A(n969), .Z(n132) );
  CTIVSVTX2 U584 ( .A(n1172), .Z(n1177) );
  B_ND2SVTX1 U585 ( .A(n1264), .B(n1263), .Z(n1265) );
  ND2SVTX6 U586 ( .A(n777), .B(n1090), .Z(n1337) );
  CTIVSVTX2 U587 ( .A(n18), .Z(n1805) );
  ND2SVTX6 U588 ( .A(n1643), .B(n827), .Z(n300) );
  NR2SVTX1 U589 ( .A(n1582), .B(n1580), .Z(n1584) );
  AO7SVTX6 U590 ( .A(n588), .B(n580), .C(n1318), .Z(n1356) );
  AO6SVTX2 U591 ( .A(n2040), .B(n2019), .C(n2018), .Z(n2020) );
  NR2SVTX6 U592 ( .A(n1630), .B(n749), .Z(n401) );
  B_ND2SVTX2 U593 ( .A(n1354), .B(n1353), .Z(n803) );
  AO6SVTX2 U594 ( .A(n2040), .B(n1372), .C(n1376), .Z(n2041) );
  NR2SVTX4 U595 ( .A(n154), .B(n917), .Z(n431) );
  AN2SVTX2 U596 ( .A(n572), .B(n1479), .Z(n570) );
  IVSVTX2 U597 ( .A(n1402), .Z(n948) );
  B_ND2SVTX2 U598 ( .A(n1982), .B(n1884), .Z(n1889) );
  CTIVSVTX4 U599 ( .A(m1[27]), .Z(n840) );
  B_ND2SVTX1 U600 ( .A(n1996), .B(n1998), .Z(n1929) );
  B_ND2SVTX2 U601 ( .A(n1982), .B(n1983), .Z(n1988) );
  IVSVTX4 U602 ( .A(n655), .Z(n1119) );
  IVSVTX0H U603 ( .A(n1783), .Z(n937) );
  ND2ASVTX6 U604 ( .A(n155), .B(n229), .Z(n655) );
  CTIVSVTX2 U605 ( .A(n1883), .Z(n1982) );
  IVSVTX2 U606 ( .A(n1723), .Z(n1812) );
  ND3SVTX4 U607 ( .A(n271), .B(n88), .C(n270), .Z(n269) );
  B_ND2SVTX2 U608 ( .A(n2051), .B(n2050), .Z(n2061) );
  IVSVTX0H U609 ( .A(n2052), .Z(n2053) );
  CTIVSVTX4 U610 ( .A(m1[1]), .Z(n155) );
  IVSVTX6 U611 ( .A(m1[1]), .Z(n939) );
  IVSVTX4 U612 ( .A(n641), .Z(n638) );
  IVSVTX6 U613 ( .A(n1915), .Z(n53) );
  B_ND2SVTX2 U614 ( .A(n1923), .B(n1922), .Z(n1925) );
  ND2SVTX6 U615 ( .A(n1716), .B(n812), .Z(m2[5]) );
  ND2SVTX6 U616 ( .A(n1847), .B(n1848), .Z(m2[9]) );
  ND2SVTX4 U617 ( .A(n987), .B(n732), .Z(n344) );
  NR2SVTX4 U618 ( .A(n1811), .B(n1826), .Z(n1848) );
  AO1SVTX4 U619 ( .A(n1670), .B(n1411), .C(n1410), .D(n1409), .Z(n1412) );
  AO17SVTX2 U620 ( .A(n991), .B(n40), .C(n990), .D(n111), .Z(n992) );
  AO3SVTX2 U621 ( .A(n1743), .B(n42), .C(n1742), .D(n1741), .Z(n1744) );
  ND2ASVTX8 U622 ( .A(n585), .B(n29), .Z(n584) );
  IVSVTX2 U623 ( .A(n1571), .Z(n1162) );
  AO6SVTX2 U624 ( .A(n1639), .B(n1640), .C(n603), .Z(n1656) );
  B_ND2SVTX2 U625 ( .A(n174), .B(n1611), .Z(n169) );
  AO2SVTX2 U626 ( .A(n1930), .B(n2036), .C(n599), .D(n816), .Z(n1950) );
  IVSVTX4 U627 ( .A(n1485), .Z(n921) );
  B_ND2SVTX2 U628 ( .A(n2071), .B(n1667), .Z(n1668) );
  ND3ABSVTX4 U629 ( .A(n494), .B(n493), .C(n492), .Z(n477) );
  ND2ASVTX4 U630 ( .A(n96), .B(n599), .Z(n279) );
  IVSVTX2 U631 ( .A(n1175), .Z(n206) );
  ND2ASVTX4 U632 ( .A(n1541), .B(n472), .Z(n1150) );
  F_ENSVTX2 U633 ( .A(n1686), .B(n1685), .Z(n1702) );
  AO7SVTX6 U634 ( .A(n984), .B(n231), .C(n983), .Z(n985) );
  IVSVTX4 U635 ( .A(n495), .Z(n492) );
  AN2SVTX4 U636 ( .A(n1170), .B(n1640), .Z(n1178) );
  IVSVTX4 U637 ( .A(n236), .Z(n238) );
  F_ENSVTX2 U638 ( .A(n1419), .B(n1415), .Z(n510) );
  IVSVTX8 U639 ( .A(n1344), .Z(n1601) );
  BFSVTX8 U640 ( .A(n287), .Z(n237) );
  CTIVSVTX6 U641 ( .A(n323), .Z(n1259) );
  ND2ASVTX4 U642 ( .A(n651), .B(n1171), .Z(n957) );
  ND3SVTX4 U643 ( .A(n632), .B(n1346), .C(n559), .Z(n389) );
  ND2ASVTX4 U644 ( .A(n1355), .B(n508), .Z(n408) );
  AO8SVTX2 U645 ( .A(n1643), .B(n1597), .C(n1870), .D(n1596), .Z(n1598) );
  IVSVTX2 U646 ( .A(n403), .Z(n1460) );
  IVSVTX4 U647 ( .A(n871), .Z(n1158) );
  B_ND2SVTX2 U648 ( .A(n1206), .B(n1205), .Z(n1208) );
  AO7SVTX6 U649 ( .A(n1218), .B(n1217), .C(n1215), .Z(n823) );
  ND2SVTX2 U650 ( .A(n1262), .B(n1261), .Z(n1256) );
  IVSVTX6 U651 ( .A(n388), .Z(n632) );
  CTIVSVTX2 U652 ( .A(n615), .Z(n1387) );
  NR2ASVTX2 U653 ( .A(n1684), .B(n1683), .Z(n1391) );
  AO7ASVTX4 U654 ( .A(n294), .B(n431), .C(n1751), .Z(n777) );
  ND2ASVTX6 U655 ( .A(n946), .B(n117), .Z(n403) );
  IVSVTX2 U656 ( .A(n688), .Z(n606) );
  NR2SVTX4 U657 ( .A(n1122), .B(n1388), .Z(n518) );
  NR2SVTX2 U658 ( .A(n182), .B(n1588), .Z(n1455) );
  B_ND2SVTX2 U659 ( .A(n1064), .B(n887), .Z(n809) );
  ND2ASVTX4 U660 ( .A(n74), .B(n1118), .Z(n615) );
  BFSVTX2 U661 ( .A(n1450), .Z(n182) );
  IVSVTX4 U662 ( .A(n1168), .Z(n47) );
  IVSVTX8 U663 ( .A(n439), .Z(n964) );
  BFSVTX2 U664 ( .A(n1382), .Z(n1684) );
  AO6SVTX4 U665 ( .A(n1804), .B(n140), .C(n858), .Z(n859) );
  B_ND2SVTX2 U666 ( .A(n1644), .B(n17), .Z(n1599) );
  AO6SVTX2 U667 ( .A(n1379), .B(n2040), .C(n1378), .Z(n1380) );
  NR2SVTX1 U668 ( .A(n1961), .B(n1708), .Z(n1712) );
  F_ND2SVTX1 U669 ( .A(n1119), .B(n1118), .Z(n705) );
  B_ND2SVTX2 U670 ( .A(n1801), .B(n140), .Z(n1809) );
  IVSVTX4 U671 ( .A(n399), .Z(n1630) );
  NR2SVTX4 U672 ( .A(n1444), .B(n1440), .Z(n1643) );
  F_AN2SVTX2 U673 ( .A(n1384), .B(n183), .Z(n1683) );
  IVSVTX10 U674 ( .A(n1131), .Z(n77) );
  NR2SVTX6 U675 ( .A(n2037), .B(n1370), .Z(n864) );
  IVSVTX6 U676 ( .A(n294), .Z(n381) );
  IVSVTX0H U677 ( .A(n1959), .Z(n1708) );
  IVSVTX0H U678 ( .A(n1367), .Z(n1690) );
  AO7SVTX4 U679 ( .A(n52), .B(n2004), .C(n272), .Z(n270) );
  CTIVSVTX2 U680 ( .A(n298), .Z(n1933) );
  CTIVSVTX2 U681 ( .A(n1703), .Z(n1967) );
  NR2SVTX4 U682 ( .A(n816), .B(n1116), .Z(n1935) );
  NR2SVTX6 U683 ( .A(n53), .B(n1916), .Z(n285) );
  IVSVTX4 U684 ( .A(n54), .Z(n113) );
  B_ND2SVTX2 U685 ( .A(n723), .B(n1897), .Z(n1680) );
  AO7SVTX4 U686 ( .A(n56), .B(n438), .C(n631), .Z(n625) );
  BFSVTX4 U687 ( .A(n1673), .Z(n1897) );
  ND3SVTX6 U688 ( .A(n1800), .B(n1799), .C(n790), .Z(m2[8]) );
  AO6SVTX2 U689 ( .A(n1745), .B(n2071), .C(n1744), .Z(n1746) );
  AO6ABSVTX4 U690 ( .A(n1902), .B(n1702), .C(n1701), .Z(n1716) );
  AO6SVTX2 U691 ( .A(n1796), .B(n2036), .C(n1795), .Z(n1797) );
  IVSVTX2 U692 ( .A(n1912), .Z(n1910) );
  NR2SVTX6 U693 ( .A(n1166), .B(n757), .Z(n1426) );
  CTIVSVTX2 U694 ( .A(n1487), .Z(n1488) );
  B_ND2SVTX2 U695 ( .A(n2022), .B(n1670), .Z(n2029) );
  B_ND2SVTX2 U696 ( .A(n1698), .B(n1670), .Z(n1699) );
  AO7NSVTX4 U697 ( .A(n1715), .B(n42), .C(n1714), .Z(n812) );
  ND2SVTX4 U698 ( .A(n1031), .B(n331), .Z(n330) );
  ND2SVTX4 U699 ( .A(n1485), .B(n1571), .Z(n471) );
  B_ND2SVTX2 U700 ( .A(n2043), .B(n1670), .Z(n2074) );
  B_ND2SVTX2 U701 ( .A(n1486), .B(n1670), .Z(n1487) );
  B_ND2SVTX2 U702 ( .A(n1943), .B(n1670), .Z(n1948) );
  AO6SVTX2 U703 ( .A(n1981), .B(n1670), .C(n1980), .Z(n1994) );
  B_ND2SVTX2 U704 ( .A(n174), .B(n1732), .Z(n1742) );
  ND3SVTX6 U705 ( .A(n35), .B(n795), .C(n1029), .Z(n333) );
  AO2SVTX2 U706 ( .A(n1533), .B(n2071), .C(n1670), .D(n1532), .Z(n1534) );
  IVSVTX6 U707 ( .A(n129), .Z(n1277) );
  B_ND2SVTX2 U708 ( .A(n1772), .B(n1670), .Z(n1800) );
  AO7SVTX2 U709 ( .A(n1408), .B(n42), .C(n1407), .Z(n1409) );
  IVSVTX2 U710 ( .A(n921), .Z(n111) );
  B_ND2SVTX2 U711 ( .A(n2071), .B(n1757), .Z(n1764) );
  IVSVTX4 U712 ( .A(n1553), .Z(n1148) );
  AO7SVTX2 U713 ( .A(n1979), .B(n60), .C(n1977), .Z(n1980) );
  B_ND2SVTX2 U714 ( .A(n2071), .B(n2027), .Z(n2028) );
  ND3ABSVTX6 U715 ( .A(n1903), .B(n494), .C(n495), .Z(n1907) );
  AO7SVTX4 U716 ( .A(n1902), .B(n510), .C(n1421), .Z(n931) );
  AO2SVTX2 U717 ( .A(n1406), .B(n2036), .C(n599), .D(n179), .Z(n1407) );
  AO2SVTX4 U718 ( .A(n498), .B(n500), .C(n390), .D(n497), .Z(n1076) );
  F_ENSVTX2 U719 ( .A(n515), .B(n876), .Z(n877) );
  B_ND2SVTX2 U720 ( .A(n1946), .B(n2071), .Z(n1947) );
  AO2SVTX2 U721 ( .A(n1514), .B(n2036), .C(n599), .D(m1[1]), .Z(n1536) );
  F_ND2SVTX1 U722 ( .A(n36), .B(n1753), .Z(n1765) );
  NR2ASVTX4 U723 ( .A(n1199), .B(n622), .Z(n621) );
  ND2SVTX4 U724 ( .A(n1342), .B(n700), .Z(n1343) );
  IVSVTX4 U725 ( .A(n1091), .Z(n59) );
  ND2ASVTX4 U726 ( .A(n708), .B(n599), .Z(n1363) );
  F_ND2SVTX1 U727 ( .A(n2048), .B(n36), .Z(n2073) );
  ND2ASVTX4 U728 ( .A(n481), .B(n599), .Z(n1421) );
  AO2SVTX2 U729 ( .A(n37), .B(n1940), .C(n174), .D(n1939), .Z(n1949) );
  IVSVTX4 U730 ( .A(n706), .Z(n494) );
  AO2SVTX2 U731 ( .A(n36), .B(n1523), .C(n174), .D(n1522), .Z(n1535) );
  ND2ASVTX4 U732 ( .A(n1000), .B(n1014), .Z(n1016) );
  IVSVTX2 U733 ( .A(n1238), .Z(n1239) );
  IVSVTX4 U734 ( .A(n714), .Z(n1001) );
  NR2ASVTX4 U735 ( .A(n672), .B(n735), .Z(n1091) );
  ND2ASVTX4 U736 ( .A(m1[23]), .B(n1055), .Z(n1054) );
  BFSVTX12 U737 ( .A(n1601), .Z(n44) );
  MUX21NSVTX4 U738 ( .A(n1339), .B(n1338), .S(n1282), .Z(n377) );
  IVSVTX4 U739 ( .A(n1259), .Z(n735) );
  IVSVTX4 U740 ( .A(n1906), .Z(n472) );
  ND3SVTX4 U741 ( .A(n842), .B(n1070), .C(n323), .Z(n1071) );
  AO7SVTX4 U742 ( .A(n1324), .B(n1323), .C(n154), .Z(n453) );
  AO6SVTX2 U743 ( .A(n1856), .B(n1684), .C(n1683), .Z(n1685) );
  ND2ASVTX6 U744 ( .A(n1000), .B(n248), .Z(n1070) );
  AO17CSVTX2 U745 ( .A(n212), .B(n1650), .C(n1649), .D(n1648), .Z(n1652) );
  B_ND2SVTX2 U746 ( .A(n1555), .B(n1565), .Z(n1903) );
  AO7CSVTX4 U747 ( .A(n730), .B(n1349), .C(n1271), .Z(n569) );
  B_ND2SVTX2 U748 ( .A(n126), .B(n1413), .Z(n1417) );
  IVSVTX2 U749 ( .A(n1541), .Z(n1542) );
  CTIVSVTX2 U750 ( .A(n1224), .Z(n1225) );
  ND2SVTX4 U751 ( .A(n1597), .B(n1870), .Z(n1650) );
  B_ND2SVTX2 U752 ( .A(n1262), .B(n1260), .Z(n1266) );
  IVSVTX4 U753 ( .A(n1049), .Z(n352) );
  ND3SVTX4 U754 ( .A(n240), .B(n106), .C(n766), .Z(n277) );
  B_ND2SVTX2 U755 ( .A(n1286), .B(n68), .Z(n1219) );
  CTIVSVTX2 U756 ( .A(n1728), .Z(n1496) );
  B_ND2SVTX2 U757 ( .A(n1462), .B(n139), .Z(n1503) );
  IVSVTX4 U758 ( .A(n1048), .Z(n351) );
  AO6SVTX6 U759 ( .A(n282), .B(n605), .C(n280), .Z(n275) );
  AO7CSVTX4 U760 ( .A(n1075), .B(n1048), .C(n99), .Z(n116) );
  B_ND2SVTX2 U761 ( .A(n826), .B(n68), .Z(n1224) );
  AO6SVTX4 U762 ( .A(n982), .B(n764), .C(n979), .Z(n763) );
  AO6SVTX6 U763 ( .A(n893), .B(n1356), .C(n892), .Z(n913) );
  IVSVTX4 U764 ( .A(n1047), .Z(n1049) );
  IVSVTX4 U765 ( .A(n1050), .Z(n63) );
  B_ND2SVTX1 U766 ( .A(n1803), .B(n409), .Z(n1807) );
  ND2SVTX4 U767 ( .A(n665), .B(n1193), .Z(n1050) );
  B_ND2SVTX2 U768 ( .A(n1169), .B(n1168), .Z(n1172) );
  ND3ABSVTX6 U769 ( .A(n928), .B(n100), .C(n460), .Z(n375) );
  B_ND2SVTX2 U770 ( .A(n1492), .B(n1491), .Z(n1500) );
  B_ND2SVTX2 U771 ( .A(n886), .B(n933), .Z(n806) );
  B_ND2SVTX2 U772 ( .A(n1061), .B(n1060), .Z(n1067) );
  AO6SVTX4 U773 ( .A(n1356), .B(n1353), .C(n1249), .Z(n579) );
  OR2SVTX2 U774 ( .A(n1333), .B(n1332), .Z(n814) );
  IVSVTX8 U775 ( .A(n506), .Z(n65) );
  IVSVTX4 U776 ( .A(n1075), .Z(n69) );
  ND2SVTX6 U777 ( .A(n74), .B(n527), .Z(n1385) );
  CTIVSVTX2 U778 ( .A(n139), .Z(n1463) );
  IVSVTX4 U779 ( .A(n1358), .Z(n73) );
  CTIVSVTX2 U780 ( .A(n1428), .Z(n1615) );
  IVSVTX4 U781 ( .A(n387), .Z(n388) );
  NR2SVTX6 U782 ( .A(n846), .B(n845), .Z(n766) );
  F_AN2SVTX2 U783 ( .A(n1643), .B(n17), .Z(n1649) );
  CTIVSVTX2 U784 ( .A(n656), .Z(n1999) );
  NR2ASVTX4 U785 ( .A(m1[24]), .B(n843), .Z(n92) );
  IVSVTX4 U786 ( .A(n1285), .Z(n68) );
  ND2SVTX6 U787 ( .A(n610), .B(n609), .Z(n949) );
  NR3SVTX6 U788 ( .A(n515), .B(n78), .C(m1[27]), .Z(n1296) );
  ND2SVTX6 U789 ( .A(n708), .B(n171), .Z(n1658) );
  IVSVTX4 U790 ( .A(n952), .Z(n1458) );
  IVSVTX2 U791 ( .A(n385), .Z(n301) );
  ND3SVTX4 U792 ( .A(n864), .B(n1372), .C(n1374), .Z(n865) );
  IVSVTX4 U793 ( .A(n1119), .Z(n74) );
  NR2SVTX6 U794 ( .A(n1957), .B(n1961), .Z(n947) );
  ND3SVTX4 U795 ( .A(n1734), .B(n463), .C(n1961), .Z(n429) );
  AO7SVTX4 U796 ( .A(n1995), .B(n1996), .C(n683), .Z(n1402) );
  B_ND2SVTX2 U797 ( .A(m1[24]), .B(m1[25]), .Z(n965) );
  B_ND2SVTX1 U798 ( .A(n1966), .B(n1965), .Z(n1974) );
  B_ND2SVTX2 U799 ( .A(n1180), .B(n1179), .Z(n807) );
  NR2SVTX4 U800 ( .A(n80), .B(n268), .Z(n267) );
  BFSVTX2 U801 ( .A(n1444), .Z(n216) );
  ND2SVTX6 U802 ( .A(n1612), .B(n1480), .Z(n563) );
  B_ND2SVTX2 U803 ( .A(n1525), .B(n1524), .Z(n1526) );
  B_ND2SVTX1 U804 ( .A(n2005), .B(n88), .Z(n1936) );
  IVSVTX2 U805 ( .A(n546), .Z(n741) );
  AO7SVTX4 U806 ( .A(n528), .B(n1518), .C(n1521), .Z(n529) );
  ND2SVTX1 U807 ( .A(n1831), .B(n1786), .Z(n1790) );
  IVSVTX10 U808 ( .A(n293), .Z(n294) );
  CTIVSVTX4 U809 ( .A(n1828), .Z(n765) );
  IVSVTX4 U810 ( .A(n527), .Z(n1118) );
  IVSVTX0H U811 ( .A(n1786), .Z(n1830) );
  CTIVSVTX2 U812 ( .A(n2024), .Z(n2055) );
  CTIVSVTX4 U813 ( .A(n1935), .Z(n88) );
  ND2ASVTX6 U814 ( .A(n297), .B(n102), .Z(n683) );
  B_ND2SVTX1 U815 ( .A(n179), .B(n1934), .Z(n2005) );
  IVSVTX4 U816 ( .A(n297), .Z(n303) );
  BFSVTX2 U817 ( .A(n1116), .Z(n179) );
  IVSVTX6 U818 ( .A(n1519), .Z(n52) );
  IVSVTX4 U819 ( .A(n218), .Z(n91) );
  ND3SVTX6 U820 ( .A(n1538), .B(n781), .C(n1154), .Z(n1366) );
  ND3SVTX4 U821 ( .A(n1540), .B(n207), .C(n558), .Z(n612) );
  NR2SVTX4 U822 ( .A(n721), .B(n530), .Z(n629) );
  CTIVSVTX2 U823 ( .A(n393), .Z(n207) );
  ND2ASVTX6 U824 ( .A(n1912), .B(n736), .Z(n1913) );
  IVSVTX2 U825 ( .A(n589), .Z(n635) );
  B_ND2SVTX2 U826 ( .A(n589), .B(n1896), .Z(n1901) );
  ND2SVTX6 U827 ( .A(n1918), .B(n1155), .Z(n1537) );
  NR2SVTX8 U828 ( .A(n1575), .B(n634), .Z(n577) );
  AO7SVTX6 U829 ( .A(n1426), .B(n1211), .C(n589), .Z(n634) );
  IVSVTX6 U830 ( .A(n249), .Z(n1151) );
  IVSVTX4 U831 ( .A(n1918), .Z(n54) );
  IVSVTX4 U832 ( .A(n1917), .Z(n55) );
  ND4ABSVTX6 U833 ( .A(n1610), .B(n170), .C(n169), .D(n168), .Z(m2[13]) );
  ND2SVTX6 U834 ( .A(n584), .B(n1210), .Z(n589) );
  IVSVTX6 U835 ( .A(n1552), .Z(n56) );
  AO6SVTX2 U836 ( .A(n1471), .B(n2071), .C(n1470), .Z(n1472) );
  AO6SVTX2 U837 ( .A(n1489), .B(n2071), .C(n1488), .Z(n1513) );
  IVSVTX2 U838 ( .A(n1609), .Z(n168) );
  NR2SVTX6 U839 ( .A(n330), .B(n332), .Z(n328) );
  ND4SVTX4 U840 ( .A(n2031), .B(n2030), .C(n2029), .D(n2028), .Z(m2[2]) );
  AO7SVTX4 U841 ( .A(n921), .B(n1162), .C(n279), .Z(n436) );
  ND4SVTX4 U842 ( .A(n2075), .B(n2074), .C(n2073), .D(n2072), .Z(m2[3]) );
  ND4SVTX4 U843 ( .A(n802), .B(n1236), .C(n1235), .D(n1234), .Z(n1244) );
  IVSVTX2 U844 ( .A(n1676), .Z(n771) );
  AO6SVTX2 U845 ( .A(n1880), .B(n1670), .C(n1879), .Z(n1894) );
  B_ND2SVTX2 U846 ( .A(n1700), .B(n1699), .Z(n1701) );
  NR3SVTX4 U847 ( .A(n1166), .B(n757), .C(n931), .Z(n932) );
  AO3ABSVTX4 U848 ( .A(n789), .B(n37), .C(n1469), .D(n1468), .Z(n1470) );
  AO7ABSVTX2 U849 ( .A(n2071), .B(n1622), .C(n1621), .Z(n170) );
  ND2SVTX6 U850 ( .A(n1363), .B(n742), .Z(n719) );
  AN2SVTX2 U851 ( .A(n1810), .B(n1670), .Z(n1811) );
  AO7SVTX4 U852 ( .A(m1[25]), .B(n670), .C(n45), .Z(n669) );
  NR2SVTX6 U853 ( .A(n295), .B(n284), .Z(n1676) );
  IVSVTX2 U854 ( .A(n1164), .Z(n496) );
  ND3SVTX4 U855 ( .A(n1362), .B(n485), .C(n487), .Z(n553) );
  IVSVTX8 U856 ( .A(n1908), .Z(n58) );
  NR2SVTX2 U857 ( .A(n1902), .B(n1512), .Z(n121) );
  IVSVTX4 U858 ( .A(n1570), .Z(n618) );
  AO6SVTX2 U859 ( .A(n1504), .B(n2036), .C(n602), .Z(n1511) );
  IVSVTX2 U860 ( .A(n456), .Z(n416) );
  ND3ASVTX6 U861 ( .A(n735), .B(n1343), .C(n176), .Z(n511) );
  IVSVTX2 U862 ( .A(n997), .Z(n457) );
  B_ND2SVTX2 U863 ( .A(n174), .B(n1774), .Z(n1799) );
  AO6SVTX2 U864 ( .A(n1875), .B(n2036), .C(n598), .Z(n1876) );
  B_ND2SVTX2 U865 ( .A(n2071), .B(n1693), .Z(n1700) );
  AO2SVTX2 U866 ( .A(n599), .B(n154), .C(n2036), .D(n1762), .Z(n1763) );
  F_ENSVTX2 U867 ( .A(n452), .B(n1749), .Z(n1766) );
  ENSVTX4 U868 ( .A(n26), .B(n411), .Z(n1274) );
  ND2SVTX4 U869 ( .A(n1033), .B(n1036), .Z(n1037) );
  F_EOSVTX2 U870 ( .A(n1844), .B(n1843), .Z(n1845) );
  AO6SVTX2 U871 ( .A(n1823), .B(n2036), .C(n601), .Z(n1824) );
  IVSVTX2 U872 ( .A(n848), .Z(n184) );
  NR2ASVTX4 U873 ( .A(m1[24]), .B(n44), .Z(n1007) );
  ND3ABSVTX6 U874 ( .A(n1078), .B(n1079), .C(n432), .Z(n1081) );
  NR3ABSVTX6 U875 ( .A(n1341), .B(n753), .C(n547), .Z(n512) );
  ND2SVTX4 U876 ( .A(n199), .B(n198), .Z(n176) );
  NR2ASVTX4 U877 ( .A(n738), .B(n44), .Z(n597) );
  F_ENSVTX2 U878 ( .A(n1466), .B(n1465), .Z(n1467) );
  ND3ASVTX6 U879 ( .A(n28), .B(n247), .C(n246), .Z(n1295) );
  IVSVTX2 U880 ( .A(n1176), .Z(n363) );
  NR3ASVTX4 U881 ( .A(n46), .B(n960), .C(n353), .Z(n962) );
  IVSVTX2 U882 ( .A(n1562), .Z(n314) );
  IVSVTX2 U883 ( .A(n1545), .Z(n101) );
  NR2SVTX6 U884 ( .A(n879), .B(n880), .Z(n915) );
  IVSVTX10 U885 ( .A(n305), .Z(n710) );
  F_EOSVTX2 U886 ( .A(n1662), .B(n1661), .Z(n1669) );
  B_ND2SVTX2 U887 ( .A(n540), .B(n1312), .Z(n1629) );
  IVSVTX2 U888 ( .A(n1070), .Z(n819) );
  AO6SVTX2 U889 ( .A(n219), .B(n1432), .C(n1431), .Z(n1433) );
  IVSVTX8 U890 ( .A(n1074), .Z(n355) );
  ND3SVTX4 U891 ( .A(n119), .B(n957), .C(n960), .Z(n958) );
  IVSVTX2 U892 ( .A(n1201), .Z(n181) );
  AO7SVTX6 U893 ( .A(n539), .B(n278), .C(n538), .Z(n97) );
  CTIVSVTX2 U894 ( .A(n1903), .Z(n493) );
  CTIVSVTX2 U895 ( .A(n1791), .Z(n1794) );
  B_ND2SVTX2 U896 ( .A(n1199), .B(n1197), .Z(n1198) );
  OR2SVTX4 U897 ( .A(n1038), .B(n1041), .Z(n1002) );
  IVSVTX2 U898 ( .A(n607), .Z(n1190) );
  CTIVSVTX6 U899 ( .A(n325), .Z(n1316) );
  NR2SVTX6 U900 ( .A(n1327), .B(n720), .Z(n538) );
  B_ND2SVTX2 U901 ( .A(n212), .B(n1650), .Z(n1507) );
  ND3SVTX4 U902 ( .A(n853), .B(n373), .C(n372), .Z(n367) );
  NR2ASVTX4 U903 ( .A(n21), .B(n1348), .Z(n1351) );
  B_ND2SVTX2 U904 ( .A(n1299), .B(n1298), .Z(n1301) );
  IVSVTX2 U905 ( .A(n116), .Z(n425) );
  ND2SVTX6 U906 ( .A(n276), .B(n277), .Z(n970) );
  AO7SVTX4 U907 ( .A(n1083), .B(n872), .C(n1085), .Z(n873) );
  B_ND2SVTX2 U908 ( .A(n1658), .B(n1305), .Z(n1662) );
  ND3ASVTX8 U909 ( .A(n686), .B(n215), .C(n214), .Z(n420) );
  NR2SVTX2 U910 ( .A(n980), .B(n979), .Z(n986) );
  IVSVTX4 U911 ( .A(n604), .Z(n276) );
  CTIVSVTX8 U912 ( .A(n1020), .Z(n61) );
  IVSVTX2 U913 ( .A(n1250), .Z(n407) );
  ND2ASVTX6 U914 ( .A(n964), .B(n369), .Z(n1298) );
  B_ND2SVTX2 U915 ( .A(n1831), .B(n1829), .Z(n1834) );
  ND2ASVTX6 U916 ( .A(n916), .B(n185), .Z(n1062) );
  NR2SVTX2 U917 ( .A(n1758), .B(n1360), .Z(n210) );
  AO7SVTX4 U918 ( .A(n677), .B(n1064), .C(n1061), .Z(n676) );
  B_ND2SVTX2 U919 ( .A(n1203), .B(n221), .Z(n1204) );
  AO6SVTX6 U920 ( .A(n679), .B(n886), .C(n678), .Z(n799) );
  AO7SVTX6 U921 ( .A(n977), .B(n1189), .C(n976), .Z(n1557) );
  NR2SVTX6 U922 ( .A(n1355), .B(n891), .Z(n911) );
  B_ND2SVTX2 U923 ( .A(n1631), .B(n399), .Z(n1638) );
  IVSVTX4 U924 ( .A(n1202), .Z(n679) );
  AO7SVTX2 U925 ( .A(n570), .B(n1615), .C(n1429), .Z(n1616) );
  NR2SVTX4 U926 ( .A(n956), .B(n1261), .Z(n1173) );
  IVSVTX2 U927 ( .A(n1215), .Z(n1216) );
  ND2ASVTX4 U928 ( .A(n1402), .B(n1401), .Z(n2033) );
  AO7ABSVTX6 U929 ( .A(n1249), .B(n718), .C(n1247), .Z(n892) );
  IVSVTX4 U930 ( .A(n854), .Z(n106) );
  IVSVTX4 U931 ( .A(n1060), .Z(n677) );
  IVSVTX4 U932 ( .A(n933), .Z(n678) );
  BFSVTX2 U933 ( .A(n1202), .Z(n221) );
  IVSVTX4 U934 ( .A(n929), .Z(n697) );
  IVSVTX4 U935 ( .A(n717), .Z(n794) );
  B_ND2SVTX2 U936 ( .A(n1506), .B(n1505), .Z(n1508) );
  ND2SVTX4 U937 ( .A(n1192), .B(n1195), .Z(n665) );
  IVSVTX4 U938 ( .A(n925), .Z(n927) );
  NR2SVTX2 U939 ( .A(n1886), .B(n1887), .Z(n1888) );
  B_ND2SVTX2 U940 ( .A(n1247), .B(n718), .Z(n1253) );
  NR2SVTX1 U941 ( .A(n1394), .B(n1395), .Z(n1398) );
  B_ND2SVTX2 U942 ( .A(n1642), .B(n1641), .Z(n1653) );
  B_ND2SVTX2 U943 ( .A(n1579), .B(n419), .Z(n1439) );
  IVSVTX4 U944 ( .A(n133), .Z(n827) );
  NR2SVTX1 U945 ( .A(n1459), .B(n1458), .Z(n1466) );
  IVSVTX4 U946 ( .A(n956), .Z(n652) );
  B_ND2SVTX2 U947 ( .A(n1429), .B(n1428), .Z(n1434) );
  CTIVSVTX2 U948 ( .A(n216), .Z(n1505) );
  IVSVTX2 U949 ( .A(n1347), .Z(n1271) );
  AO6ASVTX2 U950 ( .A(n1926), .B(n658), .C(n1119), .Z(n656) );
  AN3CSVTX6 U951 ( .A(n515), .B(n840), .C(m1[26]), .Z(n842) );
  B_ND2SVTX1 U952 ( .A(n138), .B(n14), .Z(n1607) );
  IVSVTX4 U953 ( .A(n571), .Z(n441) );
  IVSVTX4 U954 ( .A(n1317), .Z(n580) );
  AO7SVTX6 U955 ( .A(n901), .B(n1944), .C(n900), .Z(n1368) );
  F_AN2SVTX2 U956 ( .A(n1183), .B(n1184), .Z(n786) );
  CTIVSVTX2 U957 ( .A(n807), .Z(n724) );
  NR2SVTX6 U958 ( .A(n1494), .B(n1493), .Z(n290) );
  ND2SVTX6 U959 ( .A(n269), .B(n267), .Z(n1396) );
  ND3SVTX6 U960 ( .A(n941), .B(n940), .C(n942), .Z(n1401) );
  B_ND2SVTX2 U961 ( .A(n1689), .B(n1367), .Z(n1369) );
  B_ND2SVTX2 U962 ( .A(n2039), .B(n2038), .Z(n2042) );
  AO7SVTX4 U963 ( .A(n829), .B(n1777), .C(n828), .Z(n1814) );
  IVSVTX4 U964 ( .A(n1663), .Z(n686) );
  B_ND2SVTX2 U965 ( .A(n1688), .B(n51), .Z(n1692) );
  AO7SVTX4 U966 ( .A(n1506), .B(n1440), .C(n1441), .Z(n1646) );
  B_ND2SVTX1 U967 ( .A(n1872), .B(n1783), .Z(n1874) );
  F_AN2SVTX2 U968 ( .A(n1885), .B(n1982), .Z(n1886) );
  B_ND2SVTX2 U969 ( .A(n1442), .B(n1441), .Z(n1449) );
  IVSVTX0H U970 ( .A(n1719), .Z(n1476) );
  B_ND2SVTX2 U971 ( .A(n1813), .B(n1812), .Z(n1818) );
  IVSVTX2 U972 ( .A(n773), .Z(n291) );
  IVSVTX6 U973 ( .A(n563), .Z(n567) );
  B_ND2SVTX2 U974 ( .A(n414), .B(n2016), .Z(n2021) );
  B_ND2SVTX2 U975 ( .A(n1768), .B(n409), .Z(n1771) );
  B_ND2SVTX1 U976 ( .A(n2023), .B(n2054), .Z(n2026) );
  NR2SVTX1 U977 ( .A(n1932), .B(n1515), .Z(n1516) );
  B_ND2SVTX2 U978 ( .A(n2055), .B(n2052), .Z(n1945) );
  IVSVTX2 U979 ( .A(n953), .Z(n100) );
  B_ND2SVTX2 U980 ( .A(n2032), .B(n943), .Z(n2034) );
  IVSVTX4 U981 ( .A(n1110), .Z(n1107) );
  NR2SVTX1 U982 ( .A(n2053), .B(n2056), .Z(n2059) );
  NR2SVTX4 U983 ( .A(n1733), .B(n1125), .Z(n611) );
  IVSVTX2 U984 ( .A(n1813), .Z(n204) );
  IVSVTX4 U985 ( .A(n988), .Z(n78) );
  AO7SVTX4 U986 ( .A(n1959), .B(n1957), .C(n1958), .Z(n946) );
  IVSVTX10 U987 ( .A(m1[22]), .Z(n743) );
  B_ND2SVTX2 U988 ( .A(n1862), .B(n1861), .Z(n1868) );
  IVSVTX4 U989 ( .A(n1113), .Z(n681) );
  CTIVSVTX4 U990 ( .A(n1734), .Z(n81) );
  IVSVTX8 U991 ( .A(n1612), .Z(n84) );
  IVSVTX10 U992 ( .A(n1126), .Z(n85) );
  IVSVTX4 U993 ( .A(n902), .Z(n1831) );
  IVSVTX10 U994 ( .A(m1[15]), .Z(n951) );
  IVSVTX8 U995 ( .A(m1[13]), .Z(n750) );
  IVSVTX10 U996 ( .A(m1[9]), .Z(n1123) );
  IVSVTX10 U997 ( .A(m1[6]), .Z(n894) );
  IVSVTX12 U998 ( .A(n758), .Z(n759) );
  AO6ASVTX8 U999 ( .A(n1814), .B(n834), .C(n830), .Z(n1651) );
  IVSVTX8 U1000 ( .A(n758), .Z(n222) );
  ND2SVTX4 U1001 ( .A(n409), .B(n140), .Z(n867) );
  IVSVTX4 U1002 ( .A(n92), .Z(n841) );
  ND2ASVTX8 U1003 ( .A(n93), .B(n760), .Z(n843) );
  ND2SVTX4 U1004 ( .A(n94), .B(n1104), .Z(n1109) );
  ND2SVTX4 U1005 ( .A(n1116), .B(n303), .Z(n94) );
  IVSVTX2 U1006 ( .A(n95), .Z(n930) );
  AO5SVTX2 U1007 ( .A(n354), .B(m1[20]), .C(n666), .Z(n95) );
  EN3SVTX8 U1008 ( .A(m1[20]), .B(n354), .C(n96), .Z(n926) );
  ND3ASVTX6 U1009 ( .A(n1050), .B(n1046), .C(n351), .Z(n349) );
  AO7SVTX8 U1010 ( .A(n2054), .B(n2049), .C(n2051), .Z(n148) );
  CTIVSVTX4 U1011 ( .A(n453), .Z(n145) );
  AO7SVTX8 U1012 ( .A(n867), .B(n1769), .C(n859), .Z(n869) );
  AO6CSVTX8 U1013 ( .A(n39), .B(n1087), .C(n801), .Z(n1088) );
  ND4ABSVTX8 U1014 ( .A(n988), .B(n851), .C(n688), .D(n275), .Z(n607) );
  ND2SVTX4 U1015 ( .A(n716), .B(n944), .Z(n2039) );
  ND3SVTX8 U1016 ( .A(n847), .B(n896), .C(n226), .Z(n385) );
  ENSVTX8 U1017 ( .A(n786), .B(n1186), .Z(n361) );
  AO7SVTX6 U1018 ( .A(n1687), .B(n1689), .C(n1688), .Z(n1885) );
  ND2ASVTX8 U1019 ( .A(n98), .B(n1116), .Z(n1689) );
  IVSVTX4 U1020 ( .A(n944), .Z(n98) );
  ND2SVTX4 U1021 ( .A(n608), .B(n99), .Z(n707) );
  AO7CSVTX8 U1022 ( .A(n1541), .B(n811), .C(n101), .Z(n1553) );
  IVSVTX10 U1023 ( .A(n847), .Z(n666) );
  IVSVTX4 U1024 ( .A(n160), .Z(n102) );
  ND2SVTX4 U1025 ( .A(n24), .B(n103), .Z(n253) );
  ND2SVTX4 U1026 ( .A(n1401), .B(n948), .Z(n103) );
  AO6CSVTX8 U1027 ( .A(n561), .B(n55), .C(n1920), .Z(n1921) );
  IVSVTX2 U1028 ( .A(n944), .Z(n856) );
  IVSVTX4 U1029 ( .A(n104), .Z(n702) );
  ND2SVTX4 U1030 ( .A(n540), .B(n321), .Z(n104) );
  EO3SVTX8 U1031 ( .A(m1[17]), .B(n1130), .C(n354), .Z(n1142) );
  NR2SVTX2 U1032 ( .A(n605), .B(n784), .Z(n118) );
  ND2SVTX8 U1033 ( .A(n560), .B(n561), .Z(n662) );
  IVSVTX4 U1034 ( .A(n376), .Z(n105) );
  NR2SVTX4 U1035 ( .A(n105), .B(n1632), .Z(n484) );
  AO2SVTX6 U1036 ( .A(n1291), .B(n1292), .C(n800), .D(n37), .Z(n1293) );
  AO4SVTX6 U1037 ( .A(n109), .B(n195), .C(n205), .D(n107), .Z(n1423) );
  ND2ASVTX8 U1038 ( .A(n108), .B(n1178), .Z(n107) );
  NR2SVTX4 U1039 ( .A(n362), .B(n1175), .Z(n108) );
  IVSVTX4 U1040 ( .A(n1167), .Z(n109) );
  NR2SVTX8 U1041 ( .A(n539), .B(n278), .Z(n548) );
  ND2SVTX6 U1042 ( .A(n477), .B(n1163), .Z(n467) );
  CTIVSVTX12 U1043 ( .A(n817), .Z(n682) );
  AO6ABSVTX4 U1044 ( .A(n127), .B(n1022), .C(n1078), .Z(n824) );
  AO7SVTX6 U1045 ( .A(n1062), .B(n1066), .C(n799), .Z(n935) );
  ND2SVTX4 U1046 ( .A(n898), .B(n895), .Z(n684) );
  ENSVTX8 U1047 ( .A(n1925), .B(n112), .Z(m2[23]) );
  AO7SVTX8 U1048 ( .A(n1924), .B(n532), .C(n113), .Z(n112) );
  AO20SVTX8 U1049 ( .A(n147), .B(n114), .C(n146), .D(n145), .Z(n322) );
  IVSVTX4 U1050 ( .A(n1474), .Z(n890) );
  ND2SVTX2 U1051 ( .A(n1670), .B(n1620), .Z(n1621) );
  ND2SVTX6 U1052 ( .A(n1310), .B(n1311), .Z(n448) );
  ND2ASVTX8 U1053 ( .A(m1[22]), .B(n507), .Z(n575) );
  IVSVTX4 U1054 ( .A(n115), .Z(n1015) );
  ND2SVTX4 U1055 ( .A(n1013), .B(n395), .Z(n115) );
  ND2SVTX6 U1056 ( .A(n1328), .B(n1329), .Z(n147) );
  AO7SVTX4 U1057 ( .A(n1206), .B(n788), .C(n1184), .Z(n871) );
  IVSVTX4 U1058 ( .A(n1399), .Z(n156) );
  AO7SVTX6 U1059 ( .A(n1709), .B(n1710), .C(n947), .Z(n117) );
  EOSVTX8 U1060 ( .A(n986), .B(n985), .Z(n478) );
  NR2ASVTX6 U1061 ( .A(n69), .B(n1048), .Z(n348) );
  ND2SVTX4 U1062 ( .A(n1565), .B(n1554), .Z(n1541) );
  IVSVTX4 U1063 ( .A(n118), .Z(n1554) );
  NR2SVTX4 U1064 ( .A(n923), .B(n922), .Z(n977) );
  EN3SVTX8 U1065 ( .A(m1[20]), .B(n744), .C(n93), .Z(n922) );
  IVSVTX2 U1066 ( .A(n1443), .Z(n1597) );
  IVSVTX6 U1067 ( .A(n65), .Z(n427) );
  IVSVTX4 U1068 ( .A(n696), .Z(n1095) );
  EO3SVTX8 U1069 ( .A(n1123), .B(n122), .C(n860), .Z(n696) );
  ND3SVTX8 U1070 ( .A(n371), .B(n364), .C(n1302), .Z(n503) );
  ND4ABSVTX8 U1071 ( .A(n883), .B(n673), .C(n881), .D(n366), .Z(n364) );
  ND2SVTX6 U1072 ( .A(n1136), .B(n521), .Z(n1838) );
  AO6CSVTX8 U1073 ( .A(n1864), .B(n1862), .C(n1861), .Z(n1769) );
  IVSVTX4 U1074 ( .A(n1338), .Z(n123) );
  ND2ASVTX8 U1075 ( .A(n1339), .B(n123), .Z(n753) );
  IVSVTX6 U1076 ( .A(n418), .Z(n1574) );
  IVSVTX8 U1077 ( .A(n188), .Z(n1121) );
  ND3SVTX6 U1078 ( .A(n1326), .B(n1325), .C(n519), .Z(n1310) );
  IVSVTX6 U1079 ( .A(n557), .Z(n369) );
  AO4SVTX4 U1080 ( .A(n1038), .B(n1043), .C(n1042), .D(n805), .Z(n1044) );
  NR2SVTX4 U1081 ( .A(n1131), .B(n954), .Z(n916) );
  ND4SVTX4 U1082 ( .A(n1357), .B(n124), .C(n1044), .D(n1045), .Z(n331) );
  ND2SVTX4 U1083 ( .A(n125), .B(n1066), .Z(n124) );
  BFSVTX6 U1084 ( .A(n1414), .Z(n126) );
  ND3SVTX8 U1085 ( .A(n370), .B(n368), .C(n367), .Z(n371) );
  IVSVTX10 U1086 ( .A(n734), .Z(n895) );
  IVSVTX4 U1087 ( .A(n151), .Z(n130) );
  ND3SVTX6 U1088 ( .A(n130), .B(n1295), .C(n1275), .Z(n129) );
  ND2SVTX4 U1089 ( .A(n132), .B(n131), .Z(n246) );
  ND2SVTX4 U1090 ( .A(n966), .B(n967), .Z(n131) );
  ND2SVTX4 U1091 ( .A(n1642), .B(n1647), .Z(n133) );
  AO17SVTX8 U1092 ( .A(n63), .B(n1046), .C(n352), .D(n348), .Z(n1055) );
  ENSVTX8 U1093 ( .A(n1082), .B(n1081), .Z(n134) );
  AO2SVTX6 U1094 ( .A(n134), .B(n36), .C(n1076), .D(n1077), .Z(n264) );
  F_AN2SVTX2 U1095 ( .A(n1318), .B(n1317), .Z(n798) );
  ND2SVTX4 U1096 ( .A(n135), .B(n244), .Z(n1481) );
  IVSVTX4 U1097 ( .A(n759), .Z(n135) );
  AO7SVTX6 U1098 ( .A(n863), .B(n1531), .C(n1528), .Z(n1374) );
  ND2SVTX4 U1099 ( .A(n1068), .B(n917), .Z(n1215) );
  BFSVTX6 U1100 ( .A(n195), .Z(n136) );
  BFSVTX6 U1101 ( .A(n1446), .Z(n137) );
  IVSVTX4 U1102 ( .A(n1053), .Z(n746) );
  IVSVTX4 U1103 ( .A(n1240), .Z(n1242) );
  AO7CSVTX6 U1104 ( .A(n1416), .B(n1242), .C(n1241), .Z(n1243) );
  NR2SVTX4 U1105 ( .A(n1123), .B(n410), .Z(n829) );
  ENSVTX8 U1106 ( .A(n1767), .B(n780), .Z(m2[15]) );
  NR2SVTX6 U1107 ( .A(n1883), .B(n1881), .Z(n905) );
  ND2SVTX8 U1108 ( .A(n1681), .B(n1382), .Z(n188) );
  ND2SVTX6 U1109 ( .A(n261), .B(n309), .Z(n201) );
  ND3SVTX4 U1110 ( .A(n355), .B(n501), .C(m1[23]), .Z(n1059) );
  BFSVTX1 U1111 ( .A(n525), .Z(n139) );
  IVSVTX6 U1112 ( .A(n1529), .Z(n863) );
  NR2SVTX4 U1113 ( .A(n816), .B(n898), .Z(n1941) );
  ND2SVTX4 U1114 ( .A(n1384), .B(n1383), .Z(n142) );
  AO7SVTX2 U1115 ( .A(n1131), .B(n85), .C(m1[20]), .Z(n924) );
  ND2SVTX6 U1116 ( .A(n220), .B(n664), .Z(n661) );
  ND2ASVTX8 U1117 ( .A(n785), .B(n1144), .Z(n321) );
  NR4SVTX8 U1118 ( .A(n1267), .B(n144), .C(n143), .D(n1278), .Z(n1294) );
  NR2SVTX4 U1119 ( .A(n769), .B(n195), .Z(n143) );
  NR2SVTX4 U1120 ( .A(n1269), .B(n1268), .Z(n144) );
  IVSVTX12 U1121 ( .A(n733), .Z(n734) );
  AO7SVTX8 U1122 ( .A(n193), .B(n192), .C(n1345), .Z(n1127) );
  AO6SVTX8 U1123 ( .A(n899), .B(n2024), .C(n148), .Z(n900) );
  ND2SVTX4 U1124 ( .A(n620), .B(n149), .Z(n785) );
  AO7SVTX6 U1125 ( .A(n171), .B(n1345), .C(n294), .Z(n149) );
  BFSVTX1 U1126 ( .A(n1480), .Z(n150) );
  NR4ABCSVTX6 U1127 ( .A(n496), .B(n1277), .C(n1907), .D(n674), .Z(n987) );
  ND2SVTX4 U1128 ( .A(n1188), .B(n607), .Z(n151) );
  IVSVTX4 U1129 ( .A(n1413), .Z(n152) );
  AO6ASVTX8 U1130 ( .A(n152), .B(n1904), .C(n1212), .Z(n1246) );
  ND3SVTX6 U1131 ( .A(n258), .B(n1735), .C(n81), .Z(n609) );
  AO7SVTX6 U1132 ( .A(n1783), .B(n87), .C(n1781), .Z(n1735) );
  ND2SVTX4 U1133 ( .A(n1123), .B(n410), .Z(n828) );
  IVSVTX6 U1134 ( .A(n758), .Z(n259) );
  AO6SVTX6 U1135 ( .A(n241), .B(n240), .C(n821), .Z(n880) );
  NR2SVTX4 U1136 ( .A(n606), .B(n274), .Z(n1324) );
  AO1SVTX6 U1137 ( .A(n1565), .B(n1564), .C(n1563), .D(n1562), .Z(n1566) );
  ND2SVTX4 U1138 ( .A(n1304), .B(n165), .Z(n559) );
  ND2SVTX4 U1139 ( .A(n154), .B(n77), .Z(n1304) );
  NR2SVTX6 U1140 ( .A(n1576), .B(n628), .Z(n627) );
  AO6CSVTX8 U1141 ( .A(n327), .B(n540), .C(n1312), .Z(n1329) );
  ND2SVTX6 U1142 ( .A(n1111), .B(n694), .Z(n1382) );
  IVSVTX4 U1143 ( .A(n1524), .Z(n304) );
  IVSVTX8 U1144 ( .A(n889), .Z(n400) );
  NR2SVTX4 U1145 ( .A(n2032), .B(n156), .Z(n1710) );
  IVSVTX4 U1146 ( .A(n575), .Z(n157) );
  BFSVTX1 U1147 ( .A(n1802), .Z(n158) );
  ENSVTX6 U1148 ( .A(n809), .B(n935), .Z(n936) );
  NR2SVTX2 U1149 ( .A(m1[12]), .B(n889), .Z(n1444) );
  IVSVTX4 U1150 ( .A(n1768), .Z(n1804) );
  ND2SVTX4 U1151 ( .A(n1792), .B(n410), .Z(n1768) );
  NR2ASVTX2 U1152 ( .A(n1039), .B(n787), .Z(n888) );
  ND2SVTX4 U1153 ( .A(n1161), .B(n874), .Z(n1034) );
  NR2SVTX4 U1154 ( .A(n1083), .B(n1156), .Z(n874) );
  BFSVTX6 U1155 ( .A(n898), .Z(n160) );
  ND3SVTX6 U1156 ( .A(n644), .B(n643), .C(n646), .Z(n1570) );
  AO7SVTX6 U1157 ( .A(n1926), .B(n91), .C(n655), .Z(n940) );
  NR2ASVTX8 U1158 ( .A(n1676), .B(n324), .Z(n552) );
  NR2SVTX4 U1159 ( .A(n944), .B(n716), .Z(n2037) );
  BFSVTX1 U1160 ( .A(n1788), .Z(n164) );
  ND2SVTX4 U1161 ( .A(n712), .B(n72), .Z(n165) );
  AO7NSVTX4 U1162 ( .A(n1065), .B(n799), .C(n1064), .Z(n793) );
  AO7SVTX2 U1163 ( .A(n1825), .B(n1877), .C(n1824), .Z(n1826) );
  ENSVTX8 U1164 ( .A(n186), .B(n1921), .Z(m2[21]) );
  ND4ABSVTX8 U1165 ( .A(n689), .B(m1[17]), .C(n386), .D(n208), .Z(n845) );
  IVSVTX10 U1166 ( .A(m1[5]), .Z(n898) );
  IVSVTX6 U1167 ( .A(m1[18]), .Z(n293) );
  ND2SVTX4 U1168 ( .A(n25), .B(n301), .Z(n282) );
  AN2SVTX8 U1169 ( .A(n1812), .B(n1721), .Z(n834) );
  IVSVTX6 U1170 ( .A(n1123), .Z(n1775) );
  ND2SVTX4 U1171 ( .A(n259), .B(n1775), .Z(n1781) );
  ND2SVTX4 U1172 ( .A(n1126), .B(n167), .Z(n616) );
  F_AN2SVTX2 U1173 ( .A(n1085), .B(n1084), .Z(n796) );
  IVSVTX4 U1174 ( .A(n346), .Z(n211) );
  ND2ASVTX8 U1175 ( .A(n843), .B(n849), .Z(n241) );
  IVSVTX6 U1176 ( .A(n319), .Z(n1416) );
  F_ENSVTX2 U1177 ( .A(n1638), .B(n1637), .Z(n1639) );
  IVSVTX8 U1178 ( .A(n1674), .Z(n324) );
  ND2SVTX4 U1179 ( .A(n171), .B(n354), .Z(n1641) );
  ND2SVTX4 U1180 ( .A(n85), .B(n446), .Z(n1644) );
  BFSVTX1 U1181 ( .A(n1729), .Z(n172) );
  IVSVTX4 U1182 ( .A(n504), .Z(n1961) );
  ND2SVTX4 U1183 ( .A(n122), .B(n173), .Z(n504) );
  IVSVTX4 U1184 ( .A(m1[8]), .Z(n173) );
  AO6SVTX2 U1185 ( .A(n1451), .B(n1842), .C(n1452), .Z(n1454) );
  AO7ABSVTX4 U1186 ( .A(n85), .B(n211), .C(n924), .Z(n925) );
  IVSVTX4 U1187 ( .A(n1383), .Z(n694) );
  BFSVTX6 U1188 ( .A(n1917), .Z(n175) );
  IVSVTX4 U1189 ( .A(m1[12]), .Z(n713) );
  NR2ASVTX6 U1190 ( .A(n608), .B(n851), .Z(n557) );
  AO6SVTX6 U1191 ( .A(n1376), .B(n864), .C(n862), .Z(n866) );
  ND2SVTX4 U1192 ( .A(n1308), .B(n321), .Z(n452) );
  IVSVTX8 U1193 ( .A(n230), .Z(n287) );
  NR2SVTX4 U1194 ( .A(n135), .B(n860), .Z(n1777) );
  F_ND2ASVTX2 U1195 ( .A(n1388), .B(n2066), .Z(n1389) );
  ND2SVTX4 U1196 ( .A(n177), .B(n1994), .Z(m2[6]) );
  IVSVTX12 U1197 ( .A(n847), .Z(n928) );
  IVSVTX6 U1198 ( .A(n970), .Z(n1323) );
  IVSVTX4 U1199 ( .A(n792), .Z(n1114) );
  AO7ABSVTX8 U1200 ( .A(n47), .B(n994), .C(n995), .Z(n1048) );
  IVSVTX8 U1201 ( .A(m1[14]), .Z(n243) );
  AO6ASVTX8 U1202 ( .A(n1321), .B(n1320), .C(n1319), .Z(n1322) );
  ND3SVTX8 U1203 ( .A(n1551), .B(n1550), .C(n454), .Z(n394) );
  NR2SVTX4 U1204 ( .A(n1850), .B(n1849), .Z(n1851) );
  EN3SVTX8 U1205 ( .A(n758), .B(n906), .C(n860), .Z(n1850) );
  IVSVTX4 U1206 ( .A(n1272), .Z(n711) );
  NR4ABCSVTX6 U1207 ( .A(n437), .B(n1551), .C(n454), .D(n668), .Z(n631) );
  BFSVTX1 U1208 ( .A(n1383), .Z(n183) );
  ND3SVTX6 U1209 ( .A(n1142), .B(n296), .C(n321), .Z(n699) );
  IVSVTX4 U1210 ( .A(n934), .Z(n185) );
  NR2SVTX4 U1211 ( .A(n523), .B(n223), .Z(n186) );
  OR3SVTX2 U1212 ( .A(n1563), .B(n1557), .C(n1556), .Z(n791) );
  BFSVTX1 U1213 ( .A(n1627), .Z(n187) );
  IVSVTX8 U1214 ( .A(m1[18]), .Z(n708) );
  NR2SVTX4 U1215 ( .A(n1694), .B(n1951), .Z(n1863) );
  NR2ASVTX6 U1216 ( .A(n944), .B(n482), .Z(n1951) );
  IVSVTX4 U1217 ( .A(n296), .Z(n1143) );
  ND2ASVTX8 U1218 ( .A(n189), .B(n1127), .Z(n296) );
  IVSVTX4 U1219 ( .A(n1128), .Z(n189) );
  IVSVTX8 U1220 ( .A(n944), .Z(n1094) );
  AO6SVTX6 U1221 ( .A(n40), .B(n1010), .C(n534), .Z(n533) );
  BFSVTX1 U1222 ( .A(n1787), .Z(n190) );
  IVSVTX8 U1223 ( .A(n912), .Z(n227) );
  ND2SVTX4 U1224 ( .A(n1570), .B(n1163), .Z(n731) );
  AO7SVTX8 U1225 ( .A(n1758), .B(n73), .C(n1359), .Z(n1255) );
  IVSVTX8 U1226 ( .A(n77), .Z(n917) );
  AO6SVTX6 U1227 ( .A(n40), .B(n991), .C(n875), .Z(n876) );
  AO7SVTX4 U1228 ( .A(n1703), .B(n1964), .C(n1966), .Z(n836) );
  AO2ABSVTX8 U1229 ( .C(n339), .D(n340), .A(n55), .B(n1539), .Z(n338) );
  BFSVTX4 U1230 ( .A(n928), .Z(n196) );
  IVSVTX4 U1231 ( .A(n1436), .Z(n214) );
  AO6SVTX8 U1232 ( .A(n535), .B(n874), .C(n873), .Z(n1009) );
  IVSVTX4 U1233 ( .A(n197), .Z(n782) );
  ND2SVTX4 U1234 ( .A(n943), .B(n1399), .Z(n197) );
  NR2SVTX4 U1235 ( .A(n1185), .B(n788), .Z(n1161) );
  NR2SVTX4 U1236 ( .A(n76), .B(n917), .Z(n1185) );
  IVSVTX4 U1237 ( .A(n548), .Z(n198) );
  NR2SVTX4 U1238 ( .A(n753), .B(n514), .Z(n199) );
  AO7SVTX6 U1239 ( .A(n1857), .B(n1851), .C(n200), .Z(n1103) );
  AO7NSVTX4 U1240 ( .A(n34), .B(n1798), .C(n1797), .Z(n790) );
  IVSVTX2 U1241 ( .A(n1368), .Z(n1985) );
  AO7SVTX8 U1242 ( .A(n202), .B(n201), .C(n1069), .Z(n1567) );
  IVSVTX4 U1243 ( .A(n1717), .Z(n1482) );
  ND2SVTX4 U1244 ( .A(n759), .B(n675), .Z(n1717) );
  IVSVTX4 U1245 ( .A(n203), .Z(n513) );
  ND4SVTX4 U1246 ( .A(n753), .B(n1341), .C(n1340), .D(n514), .Z(n203) );
  AO3ASVTX6 U1247 ( .A(n1923), .B(n626), .C(n623), .D(n625), .Z(n630) );
  IVSVTX4 U1248 ( .A(n1004), .Z(n1005) );
  NR2ASVTX6 U1249 ( .A(n785), .B(n1144), .Z(n1145) );
  AN2SVTX8 U1250 ( .A(n1140), .B(n1139), .Z(n1588) );
  ND2SVTX4 U1251 ( .A(n1862), .B(n1863), .Z(n1802) );
  ENSVTX8 U1252 ( .A(n806), .B(n918), .Z(n1167) );
  ND2ASVTX8 U1253 ( .A(n843), .B(n849), .Z(n971) );
  ND4ABSVTX8 U1254 ( .A(n1632), .B(n385), .C(n384), .D(n383), .Z(n849) );
  ND2ASVTX8 U1255 ( .A(n347), .B(n48), .Z(n1358) );
  BFSVTX6 U1256 ( .A(n1651), .Z(n212) );
  ND3SVTX8 U1257 ( .A(n321), .B(n1141), .C(n213), .Z(n318) );
  IVSVTX4 U1258 ( .A(n509), .Z(n215) );
  IVSVTX8 U1259 ( .A(n592), .Z(n1919) );
  NR2ASVTX6 U1260 ( .A(n217), .B(n357), .Z(n1816) );
  ND2ASVTX8 U1261 ( .A(n759), .B(n860), .Z(n217) );
  ND2SVTX2 U1262 ( .A(n1654), .B(n36), .Z(n1655) );
  AO3SVTX4 U1263 ( .A(n1902), .B(n1657), .C(n1656), .D(n1655), .Z(n1671) );
  ND3ASVTX6 U1264 ( .A(n1032), .B(n334), .C(n333), .Z(n332) );
  NR3SVTX8 U1265 ( .A(n260), .B(n1537), .C(n1539), .Z(n339) );
  ND2ASVTX8 U1266 ( .A(n57), .B(n394), .Z(n1922) );
  AO7SVTX4 U1267 ( .A(m1[8]), .B(m1[10]), .C(n759), .Z(n505) );
  IVSVTX4 U1268 ( .A(n435), .Z(n1217) );
  ND2SVTX4 U1269 ( .A(n77), .B(n75), .Z(n435) );
  AN4SVTX4 U1270 ( .A(n1765), .B(n808), .C(n1764), .D(n1763), .Z(n778) );
  AO6CSVTX8 U1271 ( .A(n40), .B(n1205), .C(n1206), .Z(n1186) );
  IVSVTX4 U1272 ( .A(n1346), .Z(n730) );
  IVSVTX2 U1273 ( .A(m1[16]), .Z(n405) );
  ND2ASVTX8 U1274 ( .A(n1676), .B(n324), .Z(n551) );
  BFSVTX6 U1275 ( .A(n1430), .Z(n219) );
  NR2SVTX4 U1276 ( .A(n218), .B(n895), .Z(n1531) );
  AO7SVTX6 U1277 ( .A(n1919), .B(n1920), .C(n502), .Z(n220) );
  AO6SVTX8 U1278 ( .A(n406), .B(n404), .C(n245), .Z(n582) );
  ND2SVTX4 U1279 ( .A(n531), .B(n562), .Z(n530) );
  ND2SVTX8 U1280 ( .A(n591), .B(n361), .Z(n1420) );
  IVSVTX8 U1281 ( .A(n440), .Z(n1159) );
  ENSVTX6 U1282 ( .A(n804), .B(n250), .Z(n1754) );
  ND3SVTX8 U1283 ( .A(n1918), .B(n415), .C(n1155), .Z(n558) );
  ND2ASVTX8 U1284 ( .A(n89), .B(n400), .Z(n419) );
  NR2SVTX4 U1285 ( .A(n773), .B(n1134), .Z(n1839) );
  EN3SVTX8 U1286 ( .A(n222), .B(n1775), .C(n410), .Z(n1134) );
  ND2ASVTX8 U1287 ( .A(m1[14]), .B(n167), .Z(n1632) );
  ND2ASVTX8 U1288 ( .A(n541), .B(n1588), .Z(n1313) );
  ND2SVTX4 U1289 ( .A(n224), .B(n225), .Z(n1138) );
  EN3SVTX8 U1290 ( .A(n752), .B(m1[16]), .C(n400), .Z(n1139) );
  IVSVTX6 U1291 ( .A(n869), .Z(n565) );
  NR3ABSVTX8 U1292 ( .A(n913), .B(n914), .C(n227), .Z(n1066) );
  ND2SVTX4 U1293 ( .A(n734), .B(n898), .Z(n2054) );
  ENSVTX8 U1294 ( .A(n1427), .B(n285), .Z(m2[19]) );
  ND2SVTX4 U1295 ( .A(n1334), .B(n825), .Z(n1288) );
  ND2SVTX4 U1296 ( .A(n77), .B(n405), .Z(n1334) );
  NR4SVTX8 U1297 ( .A(n228), .B(n550), .C(n553), .D(n549), .Z(n1675) );
  NR2SVTX4 U1298 ( .A(n1361), .B(n544), .Z(n228) );
  IVSVTX4 U1299 ( .A(n297), .Z(n229) );
  AO7SVTX6 U1300 ( .A(n1446), .B(n838), .C(n1445), .Z(n235) );
  ND2SVTX8 U1301 ( .A(n287), .B(n288), .Z(n233) );
  ND2SVTX6 U1302 ( .A(n234), .B(n235), .Z(n288) );
  NR2SVTX4 U1303 ( .A(n1443), .B(n300), .Z(n234) );
  ND2SVTX4 U1304 ( .A(n1816), .B(n834), .Z(n1443) );
  IVSVTX4 U1305 ( .A(n288), .Z(n236) );
  ND2SVTX6 U1306 ( .A(n919), .B(n241), .Z(n323) );
  NR3ABSVTX8 U1307 ( .A(n1309), .B(n43), .C(n242), .Z(n449) );
  AO6SVTX1 U1308 ( .A(n1842), .B(n1311), .C(n242), .Z(n1749) );
  ND2SVTX6 U1309 ( .A(n1329), .B(n1328), .Z(n242) );
  IVSVTX12 U1310 ( .A(n243), .Z(n244) );
  IVSVTX4 U1311 ( .A(m1[14]), .Z(n675) );
  IVSVTX4 U1312 ( .A(n1978), .Z(n1640) );
  ND3SVTX4 U1313 ( .A(n1297), .B(n1978), .C(n1295), .Z(n284) );
  ND2ASVTX8 U1314 ( .A(n1257), .B(n479), .Z(n1978) );
  ND2SVTX4 U1315 ( .A(n1070), .B(n880), .Z(n1297) );
  IVSVTX4 U1316 ( .A(n971), .Z(n248) );
  AO7ABSVTX8 U1317 ( .A(n591), .B(n329), .C(n328), .Z(n249) );
  ND2ASVTX8 U1318 ( .A(n1147), .B(n249), .Z(n1918) );
  ND3ABSVTX8 U1319 ( .A(n867), .B(n1802), .C(n1696), .Z(n868) );
  ND2SVTX8 U1320 ( .A(n565), .B(n868), .Z(n1430) );
  ND2SVTX6 U1321 ( .A(n402), .B(n253), .Z(n257) );
  AO1CDSVTX8 U1322 ( .A(n257), .B(n256), .C(n397), .D(n254), .Z(n1074) );
  NR2SVTX4 U1323 ( .A(n255), .B(n745), .Z(n254) );
  NR2SVTX4 U1324 ( .A(n1602), .B(n1630), .Z(n255) );
  AO1CDSVTX8 U1325 ( .A(n1461), .B(n1501), .C(n66), .D(n401), .Z(n256) );
  ND2SVTX4 U1326 ( .A(n1124), .B(m1[8]), .Z(n1783) );
  NR2SVTX8 U1327 ( .A(n262), .B(n41), .Z(n261) );
  ND2SVTX8 U1328 ( .A(n264), .B(n263), .Z(n1165) );
  ND2SVTX8 U1329 ( .A(n591), .B(n1089), .Z(n263) );
  ND2SVTX6 U1330 ( .A(n265), .B(n537), .Z(n1575) );
  AO7SVTX8 U1331 ( .A(n1567), .B(n1165), .C(n1569), .Z(n537) );
  ND2SVTX8 U1332 ( .A(n2071), .B(n936), .Z(n1163) );
  ND2SVTX4 U1333 ( .A(n1225), .B(n232), .Z(n1230) );
  NR2SVTX8 U1334 ( .A(n90), .B(n734), .Z(n2004) );
  ND2SVTX6 U1335 ( .A(n970), .B(n607), .Z(n1344) );
  ND2SVTX4 U1336 ( .A(n70), .B(n275), .Z(n274) );
  ND2SVTX4 U1337 ( .A(n843), .B(n1000), .Z(n516) );
  ND2SVTX6 U1338 ( .A(n1326), .B(n1325), .Z(n278) );
  ND2SVTX4 U1339 ( .A(n1552), .B(n1538), .Z(n1539) );
  NR2SVTX4 U1340 ( .A(n76), .B(n281), .Z(n280) );
  NR2ASVTX6 U1341 ( .A(n376), .B(n1632), .Z(n281) );
  ND2ASVTX8 U1342 ( .A(n1747), .B(n283), .Z(n1674) );
  ND3SVTX8 U1343 ( .A(n450), .B(n322), .C(n447), .Z(n283) );
  NR2ASVTX6 U1344 ( .A(n1426), .B(n286), .Z(n1916) );
  ND2SVTX6 U1345 ( .A(n1133), .B(n1132), .Z(n1492) );
  ND2SVTX8 U1346 ( .A(n289), .B(n1315), .Z(n1452) );
  ND2SVTX8 U1347 ( .A(n1495), .B(n522), .Z(n1315) );
  NR2SVTX8 U1348 ( .A(n290), .B(n1490), .Z(n522) );
  NR2ASVTX8 U1349 ( .A(n1135), .B(n521), .Z(n1837) );
  AO7SVTX8 U1350 ( .A(n292), .B(n1490), .C(n1492), .Z(n1314) );
  NR2SVTX8 U1351 ( .A(n1133), .B(n1132), .Z(n1490) );
  AO7ABSVTX8 U1352 ( .A(n672), .B(n881), .C(n1259), .Z(n1303) );
  ND2SVTX8 U1353 ( .A(n320), .B(n1227), .Z(n1877) );
  NR2ASVTX6 U1354 ( .A(m1[5]), .B(n299), .Z(n2056) );
  NR2SVTX4 U1355 ( .A(m1[1]), .B(n299), .Z(n1926) );
  ND2SVTX4 U1356 ( .A(n342), .B(n302), .Z(n341) );
  NR2SVTX4 U1357 ( .A(n56), .B(n302), .Z(n1365) );
  AO6SVTX4 U1358 ( .A(n897), .B(n1525), .C(n304), .Z(n1944) );
  ND2SVTX4 U1359 ( .A(n939), .B(n303), .Z(n1525) );
  AO6ASVTX8 U1360 ( .A(n1002), .B(n710), .C(n1001), .Z(n306) );
  NR3ABSVTX8 U1361 ( .A(n913), .B(n914), .C(n227), .Z(n305) );
  ND3SVTX8 U1362 ( .A(n911), .B(n508), .C(n1320), .Z(n912) );
  IVSVTX12 U1363 ( .A(n894), .Z(n1106) );
  ND2SVTX4 U1364 ( .A(n905), .B(n1884), .Z(n1787) );
  ND2SVTX4 U1365 ( .A(n898), .B(n1094), .Z(n1367) );
  NR2SVTX4 U1366 ( .A(m1[8]), .B(n906), .Z(n1881) );
  NR2SVTX4 U1367 ( .A(n1123), .B(n1094), .Z(n1883) );
  AO17SVTX8 U1368 ( .A(n1063), .B(n710), .C(n310), .D(n308), .Z(n309) );
  ND2SVTX4 U1369 ( .A(n1067), .B(n793), .Z(n311) );
  ND3ABSVTX8 U1370 ( .A(n1561), .B(n314), .C(n58), .Z(n313) );
  NR3SVTX8 U1371 ( .A(n1902), .B(n1553), .C(n1566), .Z(n315) );
  NR2SVTX4 U1372 ( .A(n791), .B(n1904), .Z(n316) );
  NR2SVTX8 U1373 ( .A(n1327), .B(n318), .Z(n317) );
  ND2SVTX8 U1374 ( .A(n1729), .B(n522), .Z(n1327) );
  NR2SVTX6 U1375 ( .A(n1837), .B(n1839), .Z(n1729) );
  AO6SVTX4 U1376 ( .A(n1281), .B(n319), .C(n1280), .Z(n1292) );
  ND2SVTX6 U1377 ( .A(n1543), .B(n1544), .Z(n319) );
  IVSVTX4 U1378 ( .A(n1257), .Z(n920) );
  NR4ABCSVTX6 U1379 ( .A(n1302), .B(n1301), .C(n1303), .D(n1300), .Z(n1747) );
  ND2SVTX8 U1380 ( .A(n326), .B(n1316), .Z(n1328) );
  ND2SVTX6 U1381 ( .A(n691), .B(n1627), .Z(n325) );
  ND2SVTX6 U1382 ( .A(n289), .B(n1315), .Z(n326) );
  ND2SVTX8 U1383 ( .A(n520), .B(n1313), .Z(n327) );
  ENSVTX4 U1384 ( .A(n672), .B(n1037), .Z(n329) );
  IVSVTX4 U1385 ( .A(n561), .Z(n340) );
  ND2SVTX4 U1386 ( .A(n336), .B(n692), .Z(n337) );
  ND3SVTX4 U1387 ( .A(n1918), .B(n343), .C(n175), .Z(n342) );
  ND2SVTX6 U1388 ( .A(n345), .B(n344), .Z(n1917) );
  AO7ABSVTX2 U1389 ( .A(n2071), .B(n1167), .C(n932), .Z(n345) );
  ND2SVTX4 U1390 ( .A(n1345), .B(n211), .Z(n1359) );
  ND2SVTX4 U1391 ( .A(n350), .B(n349), .Z(n1072) );
  ND2SVTX4 U1392 ( .A(n352), .B(n351), .Z(n350) );
  IVSVTX12 U1393 ( .A(m1[11]), .Z(n758) );
  BFSVTX6 U1394 ( .A(n1074), .Z(n353) );
  ND2SVTX4 U1395 ( .A(n1012), .B(n390), .Z(n1013) );
  BFSVTX12 U1396 ( .A(m1[18]), .Z(n354) );
  ND3ABSVTX8 U1397 ( .A(n839), .B(n358), .C(n232), .Z(n1004) );
  IVSVTX12 U1398 ( .A(n1123), .Z(n1792) );
  AO7ABSVTX1 U1399 ( .A(n526), .B(n1775), .C(n728), .Z(n356) );
  NR2SVTX4 U1400 ( .A(n1423), .B(n359), .Z(n1424) );
  ND2SVTX4 U1401 ( .A(n36), .B(n360), .Z(n1422) );
  ND2SVTX4 U1402 ( .A(n726), .B(n727), .Z(n360) );
  NR2SVTX4 U1403 ( .A(n964), .B(n369), .Z(n368) );
  AO3CDSVTX8 U1404 ( .A(n65), .B(n375), .C(n988), .D(n556), .Z(n370) );
  ND2ASVTX8 U1405 ( .A(n76), .B(n374), .Z(n373) );
  IVSVTX4 U1406 ( .A(n766), .Z(n374) );
  NR3ABSVTX8 U1407 ( .A(n376), .B(n463), .C(n382), .Z(n384) );
  NR3SVTX8 U1408 ( .A(n738), .B(m1[10]), .C(n835), .Z(n376) );
  ND2SVTX4 U1409 ( .A(n377), .B(n43), .Z(n1280) );
  ND2SVTX4 U1410 ( .A(n491), .B(n378), .Z(n1282) );
  IVSVTX4 U1411 ( .A(n1279), .Z(n378) );
  NR2ASVTX8 U1412 ( .A(n1141), .B(n1450), .Z(n1627) );
  NR2SVTX8 U1413 ( .A(n1140), .B(n1139), .Z(n1450) );
  ND3SVTX8 U1414 ( .A(n1506), .B(n1462), .C(n1129), .Z(n1140) );
  NR2SVTX4 U1415 ( .A(n380), .B(n1142), .Z(n747) );
  ND2SVTX4 U1416 ( .A(n1128), .B(n1127), .Z(n380) );
  ND2SVTX4 U1417 ( .A(n77), .B(n381), .Z(n382) );
  IVSVTX4 U1418 ( .A(n845), .Z(n383) );
  ND2SVTX6 U1419 ( .A(n928), .B(n633), .Z(n387) );
  IVSVTX4 U1420 ( .A(n1074), .Z(n390) );
  NR2ASVTX6 U1421 ( .A(n1759), .B(n1074), .Z(n391) );
  ND2ASVTX8 U1422 ( .A(n57), .B(n394), .Z(n1155) );
  ND2SVTX4 U1423 ( .A(n455), .B(n394), .Z(n393) );
  NR2SVTX4 U1424 ( .A(m1[24]), .B(n1014), .Z(n395) );
  NR2SVTX4 U1425 ( .A(n60), .B(n396), .Z(n1017) );
  NR2SVTX4 U1426 ( .A(n1000), .B(n1013), .Z(n396) );
  ND2SVTX4 U1427 ( .A(n1457), .B(n1458), .Z(n398) );
  ND2SVTX4 U1428 ( .A(n952), .B(n525), .Z(n739) );
  IVSVTX4 U1429 ( .A(n419), .Z(n404) );
  ND2SVTX6 U1430 ( .A(n1579), .B(n406), .Z(n509) );
  ND2SVTX2 U1431 ( .A(n1578), .B(n406), .Z(n1586) );
  ND2SVTX4 U1432 ( .A(n407), .B(n508), .Z(n768) );
  AO7SVTX6 U1433 ( .A(n408), .B(n1248), .C(n704), .Z(n703) );
  ND2SVTX4 U1434 ( .A(n1123), .B(m1[12]), .Z(n409) );
  AO6SVTX4 U1435 ( .A(n1430), .B(n1273), .C(n412), .Z(n411) );
  AO7SVTX6 U1436 ( .A(n413), .B(n64), .C(n568), .Z(n412) );
  IVSVTX4 U1437 ( .A(n711), .Z(n413) );
  ND2SVTX4 U1438 ( .A(n273), .B(n299), .Z(n414) );
  ND2SVTX8 U1439 ( .A(n441), .B(n442), .Z(n1659) );
  AO7ABSVTX6 U1440 ( .A(n613), .B(n1568), .C(n418), .Z(n415) );
  ND3ABSVTX8 U1441 ( .A(n1153), .B(n1152), .C(n1151), .Z(n418) );
  ND3ABSVTX8 U1442 ( .A(n997), .B(n416), .C(n417), .Z(n455) );
  ND2SVTX4 U1443 ( .A(n481), .B(n48), .Z(n825) );
  IVSVTX4 U1444 ( .A(n690), .Z(n417) );
  ND2ASVTX8 U1445 ( .A(n195), .B(n1003), .Z(n1551) );
  ND2SVTX4 U1446 ( .A(n1918), .B(n418), .Z(n663) );
  NR2SVTX4 U1447 ( .A(n686), .B(n582), .Z(n422) );
  NR2SVTX4 U1448 ( .A(n685), .B(n422), .Z(n421) );
  NR2SVTX8 U1449 ( .A(n890), .B(n687), .Z(n1436) );
  ND2SVTX6 U1450 ( .A(n652), .B(n1255), .Z(n1046) );
  F_IVSVTX1 U1451 ( .A(m1[16]), .Z(n423) );
  ND2SVTX4 U1452 ( .A(n996), .B(n1171), .Z(n424) );
  ND2SVTX6 U1453 ( .A(n590), .B(n426), .Z(n642) );
  ND4ABSVTX8 U1454 ( .A(n851), .B(n968), .C(n427), .D(n818), .Z(n878) );
  NR3ABSVTX8 U1455 ( .A(n461), .B(n428), .C(n429), .Z(n506) );
  ND3SVTX4 U1456 ( .A(n1233), .B(n1232), .C(n320), .Z(n1234) );
  AO6SVTX8 U1457 ( .A(n1969), .B(n837), .C(n836), .Z(n1445) );
  ND3SVTX8 U1458 ( .A(n32), .B(n669), .C(n490), .Z(n690) );
  IVSVTX12 U1459 ( .A(m1[10]), .Z(n906) );
  ND2SVTX4 U1460 ( .A(n12), .B(m1[16]), .Z(n1441) );
  ND2SVTX4 U1461 ( .A(n405), .B(n86), .Z(n1317) );
  ND2SVTX4 U1462 ( .A(m1[16]), .B(n244), .Z(n1128) );
  ND2SVTX4 U1463 ( .A(n193), .B(n1131), .Z(n1751) );
  ND2SVTX4 U1464 ( .A(n433), .B(n233), .Z(n432) );
  ND2ASVTX8 U1465 ( .A(n1021), .B(n61), .Z(n1080) );
  ND2ASVTX8 U1466 ( .A(n434), .B(n826), .Z(n1020) );
  NR2ASVTX6 U1467 ( .A(n1025), .B(n1181), .Z(n1079) );
  AO6ASVTX8 U1468 ( .A(n434), .B(n1286), .C(n823), .Z(n1181) );
  ND2SVTX4 U1469 ( .A(n68), .B(n435), .Z(n434) );
  IVSVTX4 U1470 ( .A(n631), .Z(n1923) );
  IVSVTX4 U1471 ( .A(n455), .Z(n438) );
  ND2SVTX4 U1472 ( .A(n988), .B(n608), .Z(n439) );
  AO7SVTX8 U1473 ( .A(n1160), .B(n1159), .C(n31), .Z(n1207) );
  ND3SVTX8 U1474 ( .A(n565), .B(n64), .C(n868), .Z(n440) );
  AO3SVTX6 U1475 ( .A(n1659), .B(n1660), .C(n30), .D(n21), .Z(n1160) );
  AO17SVTX8 U1476 ( .A(n1482), .B(n567), .C(n566), .D(n1428), .Z(n442) );
  NR2SVTX4 U1477 ( .A(n1614), .B(n443), .Z(n1660) );
  ND2SVTX4 U1478 ( .A(n444), .B(n1428), .Z(n443) );
  IVSVTX4 U1479 ( .A(n1537), .Z(n576) );
  NR2SVTX4 U1480 ( .A(n1719), .B(n445), .Z(n687) );
  IVSVTX4 U1481 ( .A(n1475), .Z(n445) );
  ND2ASVTX8 U1482 ( .A(m1[12]), .B(n446), .Z(n1475) );
  ENSVTX8 U1483 ( .A(n798), .B(n1322), .Z(n1756) );
  ND2SVTX4 U1484 ( .A(n1754), .B(n503), .Z(n450) );
  ND2SVTX8 U1485 ( .A(n919), .B(n971), .Z(n479) );
  ND2SVTX4 U1486 ( .A(n1552), .B(n455), .Z(n1577) );
  ND2SVTX4 U1487 ( .A(n2036), .B(n998), .Z(n456) );
  ND2ASVTX8 U1488 ( .A(n457), .B(n690), .Z(n1552) );
  ND4ABCSVTX8 U1489 ( .A(m1[27]), .B(m1[24]), .C(n883), .D(n971), .Z(n884) );
  IVSVTX4 U1490 ( .A(n882), .Z(n883) );
  NR2ASVTX6 U1491 ( .A(m1[26]), .B(n515), .Z(n882) );
  IVSVTX4 U1492 ( .A(n1188), .Z(n1330) );
  ND2SVTX4 U1493 ( .A(n710), .B(n888), .Z(n458) );
  ND2SVTX4 U1494 ( .A(n459), .B(n715), .Z(n835) );
  IVSVTX4 U1495 ( .A(m1[7]), .Z(n459) );
  NR4SVTX8 U1496 ( .A(n752), .B(n1519), .C(n816), .D(n889), .Z(n461) );
  ND2SVTX6 U1497 ( .A(n1214), .B(n1213), .Z(n755) );
  ND2SVTX8 U1498 ( .A(n335), .B(n465), .Z(n1214) );
  ENSVTX8 U1499 ( .A(n1204), .B(n710), .Z(n465) );
  ND2SVTX6 U1500 ( .A(n469), .B(n466), .Z(n1911) );
  NR3SVTX8 U1501 ( .A(n618), .B(n468), .C(n467), .Z(n466) );
  IVSVTX4 U1502 ( .A(n470), .Z(n469) );
  ND2SVTX4 U1503 ( .A(n474), .B(n477), .Z(n674) );
  IVSVTX4 U1504 ( .A(n480), .Z(n974) );
  ND2SVTX4 U1505 ( .A(n480), .B(n972), .Z(n1565) );
  AO5ASVTX8 U1506 ( .B(n605), .A(n481), .C(n83), .Z(n480) );
  ND2SVTX8 U1507 ( .A(n708), .B(n226), .Z(n1194) );
  ND3SVTX8 U1508 ( .A(n484), .B(n49), .C(n507), .Z(n854) );
  ND2SVTX4 U1509 ( .A(n1357), .B(n486), .Z(n485) );
  F_ENSVTX2 U1510 ( .A(n803), .B(n703), .Z(n486) );
  F_EOSVTX2 U1511 ( .A(n1352), .B(n489), .Z(n488) );
  ND2SVTX4 U1512 ( .A(n591), .B(n877), .Z(n490) );
  ND2SVTX6 U1513 ( .A(n1004), .B(n671), .Z(n670) );
  AO7SVTX8 U1514 ( .A(n1337), .B(n1279), .C(n491), .Z(n1556) );
  IVSVTX4 U1515 ( .A(n811), .Z(n1564) );
  NR2SVTX4 U1516 ( .A(n69), .B(n499), .Z(n498) );
  ND2SVTX4 U1517 ( .A(n501), .B(n355), .Z(n500) );
  IVSVTX4 U1518 ( .A(n746), .Z(n501) );
  IVSVTX4 U1519 ( .A(n523), .Z(n502) );
  ND2SVTX4 U1520 ( .A(n1106), .B(n307), .Z(n1101) );
  ND2SVTX4 U1521 ( .A(n1116), .B(n307), .Z(n1393) );
  ND2ASVTX8 U1522 ( .A(m1[8]), .B(n90), .Z(n1688) );
  IVSVTX12 U1523 ( .A(n750), .Z(n752) );
  EN3SVTX8 U1524 ( .A(m1[16]), .B(n1131), .C(n294), .Z(n1144) );
  AO7SVTX6 U1525 ( .A(n509), .B(n1436), .C(n582), .Z(n517) );
  AO6CSVTX8 U1526 ( .A(n1556), .B(n126), .C(n1189), .Z(n1415) );
  IVSVTX4 U1527 ( .A(n548), .Z(n1842) );
  NR3SVTX8 U1528 ( .A(n512), .B(n513), .C(n511), .Z(n549) );
  ND2SVTX4 U1529 ( .A(n1296), .B(n516), .Z(n604) );
  AO6SVTX4 U1530 ( .A(n517), .B(n67), .C(n1356), .Z(n704) );
  AO6SVTX1 U1531 ( .A(n1435), .B(n508), .C(n517), .Z(n1665) );
  ND3SVTX8 U1532 ( .A(n1120), .B(n518), .C(n1121), .Z(n519) );
  ND2SVTX6 U1533 ( .A(n1099), .B(n1098), .Z(n1849) );
  EN3SVTX8 U1534 ( .A(m1[10]), .B(n1123), .C(n1102), .Z(n1853) );
  ND2SVTX4 U1535 ( .A(n1101), .B(n1100), .Z(n1854) );
  ND2SVTX4 U1536 ( .A(n2011), .B(n1115), .Z(n1388) );
  EO3SVTX8 U1537 ( .A(n1124), .B(n89), .C(n713), .Z(n521) );
  EO3SVTX8 U1538 ( .A(n1130), .B(n564), .C(n82), .Z(n1132) );
  EN3SVTX8 U1539 ( .A(m1[14]), .B(m1[17]), .C(m1[16]), .Z(n619) );
  IVSVTX2 U1540 ( .A(n537), .Z(n523) );
  ND2SVTX4 U1541 ( .A(n82), .B(n713), .Z(n525) );
  ND2SVTX4 U1542 ( .A(n1457), .B(n1462), .Z(n524) );
  ND2SVTX8 U1543 ( .A(n244), .B(n526), .Z(n1462) );
  ENSVTX8 U1544 ( .A(m1[1]), .B(n895), .Z(n1518) );
  EN3SVTX8 U1545 ( .A(n716), .B(n1934), .C(n1116), .Z(n527) );
  ND2SVTX4 U1546 ( .A(n1385), .B(n1938), .Z(n614) );
  ND2SVTX4 U1547 ( .A(n1517), .B(n529), .Z(n1938) );
  ND2SVTX4 U1548 ( .A(n528), .B(n1518), .Z(n1517) );
  NR2SVTX4 U1549 ( .A(n631), .B(n1577), .Z(n531) );
  IVSVTX8 U1550 ( .A(n562), .Z(n532) );
  IVSVTX4 U1551 ( .A(n559), .Z(n1349) );
  NR2SVTX4 U1552 ( .A(n672), .B(n1009), .Z(n534) );
  IVSVTX4 U1553 ( .A(n1158), .Z(n535) );
  ND2SVTX4 U1554 ( .A(n1254), .B(n536), .Z(n1197) );
  NR2SVTX4 U1555 ( .A(n981), .B(n980), .Z(n1025) );
  NR2SVTX4 U1556 ( .A(m1[20]), .B(m1[23]), .Z(n981) );
  ND2SVTX4 U1557 ( .A(n748), .B(n1143), .Z(n540) );
  IVSVTX4 U1558 ( .A(n1587), .Z(n542) );
  ND2ASVTX8 U1559 ( .A(n71), .B(n1137), .Z(n1587) );
  AO7SVTX4 U1560 ( .A(n462), .B(n526), .C(n12), .Z(n543) );
  NR2SVTX4 U1561 ( .A(n752), .B(m1[16]), .Z(n1440) );
  ND2SVTX4 U1562 ( .A(n752), .B(n462), .Z(n1813) );
  ND2SVTX4 U1563 ( .A(n12), .B(n889), .Z(n1457) );
  ND2SVTX4 U1564 ( .A(n1340), .B(n548), .Z(n547) );
  AO3SVTX6 U1565 ( .A(n1675), .B(n552), .C(n551), .D(n1672), .Z(n555) );
  ND3SVTX8 U1566 ( .A(n1673), .B(n1896), .C(n555), .Z(n587) );
  ND2SVTX6 U1567 ( .A(n1293), .B(n1294), .Z(n1673) );
  ND2ASVTX8 U1568 ( .A(n634), .B(n587), .Z(n561) );
  AO6SVTX8 U1569 ( .A(n1556), .B(n62), .C(n1557), .Z(n811) );
  NR2ASVTX6 U1570 ( .A(n775), .B(n850), .Z(n818) );
  ND2SVTX8 U1571 ( .A(n577), .B(n587), .Z(n562) );
  ND2ASVTX8 U1572 ( .A(n951), .B(n564), .Z(n1480) );
  IVSVTX12 U1573 ( .A(m1[12]), .Z(n564) );
  ND2SVTX4 U1574 ( .A(m1[12]), .B(n855), .Z(n1479) );
  AO7SVTX6 U1575 ( .A(n1429), .B(n84), .C(n1613), .Z(n571) );
  NR2ASVTX6 U1576 ( .A(m1[27]), .B(n878), .Z(n879) );
  ND2SVTX4 U1577 ( .A(n574), .B(n1556), .Z(n1221) );
  IVSVTX4 U1578 ( .A(n574), .Z(n1237) );
  ND2SVTX4 U1579 ( .A(n1353), .B(n718), .Z(n891) );
  ND2SVTX4 U1580 ( .A(n1353), .B(n67), .Z(n1250) );
  ND2SVTX4 U1581 ( .A(n211), .B(n48), .Z(n1353) );
  NR3SVTX8 U1582 ( .A(n584), .B(n1246), .C(n755), .Z(n583) );
  ND3SVTX8 U1583 ( .A(n654), .B(n895), .C(n675), .Z(n586) );
  MUX21NSVTX2 U1584 ( .A(n1266), .B(n1265), .S(n355), .Z(n1268) );
  ND2SVTX4 U1585 ( .A(n171), .B(n709), .Z(n588) );
  NR3SVTX4 U1586 ( .A(m1[24]), .B(m1[27]), .C(n850), .Z(n590) );
  NR3ABSVTX8 U1587 ( .A(n593), .B(n664), .C(n662), .Z(n659) );
  IVSVTX4 U1588 ( .A(n223), .Z(n593) );
  IVSVTX4 U1589 ( .A(n594), .Z(n1069) );
  NR2ASVTX6 U1590 ( .A(n1068), .B(n44), .Z(n594) );
  NR2ASVTX6 U1591 ( .A(n1792), .B(n44), .Z(n595) );
  NR2SVTX4 U1592 ( .A(n741), .B(n611), .Z(n610) );
  ND2SVTX4 U1593 ( .A(m1[12]), .B(n462), .Z(n1125) );
  ND2SVTX4 U1594 ( .A(n615), .B(n614), .Z(n1120) );
  ND2SVTX4 U1595 ( .A(n218), .B(m1[2]), .Z(n1927) );
  ND2ASVTX8 U1596 ( .A(n347), .B(n954), .Z(n1192) );
  ND2SVTX4 U1597 ( .A(n1345), .B(n171), .Z(n620) );
  IVSVTX4 U1598 ( .A(n1922), .Z(n624) );
  NR3SVTX8 U1599 ( .A(n630), .B(n629), .C(n627), .Z(m2[24]) );
  IVSVTX4 U1600 ( .A(n354), .Z(n633) );
  IVSVTX6 U1601 ( .A(n640), .Z(n1427) );
  MUX21NSVTX6 U1602 ( .A(n1916), .B(n53), .S(n641), .Z(n636) );
  ND3SVTX4 U1603 ( .A(n1427), .B(n1915), .C(n638), .Z(n637) );
  ND2SVTX4 U1604 ( .A(n645), .B(n955), .Z(n644) );
  NR2SVTX4 U1605 ( .A(n60), .B(n962), .Z(n646) );
  NR2SVTX4 U1606 ( .A(n650), .B(n648), .Z(n647) );
  IVSVTX4 U1607 ( .A(n1161), .Z(n649) );
  AO7SVTX6 U1608 ( .A(n649), .B(n31), .C(n1158), .Z(n650) );
  ND3SVTX6 U1609 ( .A(n1302), .B(n364), .C(n371), .Z(n1485) );
  ND2SVTX2 U1610 ( .A(n653), .B(n1695), .Z(n1697) );
  IVSVTX4 U1611 ( .A(n663), .Z(n664) );
  AO7ABSVTX4 U1612 ( .A(n223), .B(n663), .C(n661), .Z(n660) );
  ND2ASVTX8 U1613 ( .A(n1910), .B(n1911), .Z(n1920) );
  IVSVTX4 U1614 ( .A(n1254), .Z(n1195) );
  ND2SVTX4 U1615 ( .A(n1254), .B(n1194), .Z(n1262) );
  ND2ASVTX8 U1616 ( .A(n708), .B(n79), .Z(n1254) );
  ND2SVTX8 U1617 ( .A(n515), .B(n1000), .Z(n851) );
  ND2SVTX4 U1618 ( .A(n691), .B(n1627), .Z(n720) );
  ND2ASVTX8 U1619 ( .A(n928), .B(n917), .Z(n1202) );
  NR2ASVTX6 U1620 ( .A(m1[24]), .B(n670), .Z(n1008) );
  IVSVTX4 U1621 ( .A(n1006), .Z(n671) );
  ND2ASVTX8 U1622 ( .A(n75), .B(n849), .Z(n881) );
  AO7ABSVTX8 U1623 ( .A(n672), .B(n881), .C(n885), .Z(n1188) );
  ND2SVTX4 U1624 ( .A(n1000), .B(n853), .Z(n673) );
  IVSVTX6 U1625 ( .A(m1[26]), .Z(n988) );
  ND2SVTX4 U1626 ( .A(n196), .B(n556), .Z(n1064) );
  IVSVTX4 U1627 ( .A(n886), .Z(n934) );
  AO6ABSVTX6 U1628 ( .A(n680), .B(n799), .C(n676), .Z(n1040) );
  ND2ASVTX6 U1629 ( .A(n928), .B(n83), .Z(n887) );
  ND2SVTX4 U1630 ( .A(n792), .B(n681), .Z(n2010) );
  IVSVTX4 U1631 ( .A(n684), .Z(n1995) );
  AO6SVTX4 U1632 ( .A(n845), .B(n1068), .C(n707), .Z(n688) );
  ND2SVTX4 U1633 ( .A(n938), .B(n951), .Z(n689) );
  IVSVTX4 U1634 ( .A(n747), .Z(n691) );
  NR2SVTX6 U1635 ( .A(n1365), .B(n1366), .Z(m2[26]) );
  ND2SVTX6 U1636 ( .A(n1552), .B(n692), .Z(n1154) );
  AO6SVTX8 U1637 ( .A(n1855), .B(n1112), .C(n1103), .Z(n1326) );
  ND2SVTX1 U1638 ( .A(n693), .B(n1882), .Z(n1891) );
  ND2SVTX8 U1639 ( .A(n975), .B(n1414), .Z(n1558) );
  ND2ASVTX8 U1640 ( .A(n930), .B(n697), .Z(n1414) );
  ND2ASVTX8 U1641 ( .A(n923), .B(n698), .Z(n975) );
  IVSVTX4 U1642 ( .A(n922), .Z(n698) );
  ND2ASVTX8 U1643 ( .A(n1145), .B(n699), .Z(n701) );
  ND2SVTX6 U1644 ( .A(n1341), .B(n1340), .Z(n700) );
  ND2SVTX8 U1645 ( .A(n1452), .B(n1336), .Z(n1341) );
  AO6SVTX8 U1646 ( .A(n702), .B(n1623), .C(n701), .Z(n1340) );
  ND2SVTX4 U1647 ( .A(n1035), .B(n39), .Z(n1036) );
  AO8ASVTX2 U1648 ( .A(n1737), .B(n81), .C(n1873), .D(n1736), .Z(n1738) );
  AO7SVTX2 U1649 ( .A(n1323), .B(n1190), .C(n917), .Z(n1191) );
  AO7SVTX4 U1650 ( .A(n1303), .B(n1221), .C(n1191), .Z(n1241) );
  EN3SVTX8 U1651 ( .A(n715), .B(n1106), .C(n1105), .Z(n1110) );
  F_ND2SVTX0H U1652 ( .A(n1519), .B(m1[1]), .Z(n1931) );
  ND2SVTX2 U1653 ( .A(n259), .B(n244), .Z(n1722) );
  NR2SVTX2 U1654 ( .A(m1[10]), .B(n938), .Z(n857) );
  AO7SVTX6 U1655 ( .A(n1751), .B(n1332), .C(n1331), .Z(n1286) );
  AO7ABSVTX4 U1656 ( .A(n21), .B(n1659), .C(n1349), .Z(n1350) );
  IVSVTX10 U1657 ( .A(m1[21]), .Z(n847) );
  AO2SVTX2 U1658 ( .A(n820), .B(m1[27]), .C(n819), .D(n783), .Z(n822) );
  OR2ABSVTX8 U1659 ( .A(n1188), .B(n915), .Z(n2071) );
  F_IVSVTX0H U1660 ( .A(n2010), .Z(n2064) );
  AO7SVTX2 U1661 ( .A(n1961), .B(n1960), .C(n1959), .Z(n1962) );
  ND2SVTX4 U1662 ( .A(n1123), .B(n1094), .Z(n1983) );
  F_ND2ASVTX2 U1663 ( .A(m1[4]), .B(m1[1]), .Z(n1528) );
  IVSVTX2 U1664 ( .A(n1025), .Z(n1021) );
  ND2SVTX4 U1665 ( .A(n1345), .B(n77), .Z(n1354) );
  IVSVTX4 U1666 ( .A(n1354), .Z(n1249) );
  F_ND2SVTX0H U1667 ( .A(n1347), .B(n1346), .Z(n1352) );
  IVSVTX4 U1668 ( .A(n1916), .Z(n1914) );
  EOSVTX4 U1669 ( .A(n1419), .B(n1418), .Z(n1425) );
  ND2ASVTX8 U1670 ( .A(n953), .B(n708), .Z(n718) );
  IVSVTX2 U1671 ( .A(m1[21]), .Z(n954) );
  AO7SVTX8 U1672 ( .A(n767), .B(n768), .C(n1251), .Z(n1252) );
  NR2SVTX2 U1673 ( .A(m1[8]), .B(n682), .Z(n1395) );
  ND3ABSVTX8 U1674 ( .A(n1919), .B(n1574), .C(n1573), .Z(n721) );
  ND3SVTX8 U1675 ( .A(n1572), .B(n1909), .C(n1917), .Z(n1573) );
  NR2ASVTX6 U1676 ( .A(n1357), .B(n769), .Z(n722) );
  AO7SVTX2 U1677 ( .A(n722), .B(n719), .C(n1364), .Z(n723) );
  ND2SVTX2 U1678 ( .A(n807), .B(n1182), .Z(n726) );
  ND2SVTX4 U1679 ( .A(n724), .B(n725), .Z(n727) );
  IVSVTX2 U1680 ( .A(n1182), .Z(n725) );
  AO7SVTX2 U1681 ( .A(n1776), .B(n1778), .C(n1869), .Z(n1779) );
  ND2SVTX4 U1682 ( .A(n83), .B(n196), .Z(n995) );
  ND2ASVTX8 U1683 ( .A(n953), .B(n744), .Z(n1168) );
  AO7SVTX4 U1684 ( .A(n1417), .B(n1908), .C(n1415), .Z(n1418) );
  AO4SVTX2 U1685 ( .A(n811), .B(n1546), .C(n672), .D(n1545), .Z(n1547) );
  ND2SVTX4 U1686 ( .A(n742), .B(n1277), .Z(n1278) );
  ENSVTX8 U1687 ( .A(n796), .B(n1088), .Z(n1089) );
  AO7SVTX4 U1688 ( .A(n839), .B(n166), .C(n824), .Z(n1006) );
  ND2SVTX2 U1689 ( .A(n244), .B(m1[16]), .Z(n1602) );
  ND2SVTX4 U1690 ( .A(n761), .B(m1[20]), .Z(n933) );
  AO7SVTX2 U1691 ( .A(n1082), .B(n1078), .C(m1[23]), .Z(n1026) );
  IVSVTX4 U1692 ( .A(n1911), .Z(n736) );
  NR2SVTX2 U1693 ( .A(n738), .B(n1775), .Z(n737) );
  NR2SVTX2 U1694 ( .A(n738), .B(n1775), .Z(n1972) );
  IVSVTX4 U1695 ( .A(n825), .Z(n1332) );
  ND2SVTX4 U1696 ( .A(n1831), .B(n1828), .Z(n909) );
  NR2SVTX4 U1697 ( .A(n909), .B(n1787), .Z(n903) );
  NR2SVTX2 U1698 ( .A(n218), .B(m1[2]), .Z(n1117) );
  ND3SVTX2 U1699 ( .A(m1[23]), .B(n61), .C(n1025), .Z(n1028) );
  IVSVTX4 U1700 ( .A(n1435), .Z(n767) );
  ND2SVTX2 U1701 ( .A(n1105), .B(n1775), .Z(n1099) );
  ND3ABSVTX4 U1702 ( .A(n1283), .B(n1339), .C(n1416), .Z(n1291) );
  NR2SVTX2 U1703 ( .A(m1[10]), .B(m1[8]), .Z(n1782) );
  CTIVSVTX4 U1704 ( .A(n1554), .Z(n1561) );
  IVSVTX2 U1705 ( .A(n1135), .Z(n1136) );
  NR2SVTX2 U1706 ( .A(n1782), .B(n87), .Z(n1820) );
  ND2SVTX2 U1707 ( .A(n840), .B(n882), .Z(n821) );
  AO7ABSVTX4 U1708 ( .A(n2033), .B(n24), .C(n1460), .Z(n1873) );
  IVSVTX2 U1709 ( .A(n1565), .Z(n1560) );
  NR2SVTX2 U1710 ( .A(n672), .B(n1034), .Z(n1010) );
  NR2SVTX2 U1711 ( .A(n1760), .B(n545), .Z(n1761) );
  IVSVTX4 U1712 ( .A(n1642), .Z(n831) );
  F_ND2ASVTX2 U1713 ( .A(n1284), .B(n1219), .Z(n1228) );
  IVSVTX2 U1714 ( .A(n1218), .Z(n1284) );
  F_ND2ASVTX2 U1715 ( .A(n672), .B(n1079), .Z(n1027) );
  AO6SVTX2 U1716 ( .A(n1856), .B(n1121), .C(n1855), .Z(n1990) );
  AO6SVTX1 U1717 ( .A(n1873), .B(n1820), .C(n1735), .Z(n1821) );
  NR2SVTX0H U1718 ( .A(n741), .B(n1733), .Z(n1739) );
  ND2SVTX4 U1719 ( .A(n1126), .B(n244), .Z(n1613) );
  ND2SVTX4 U1720 ( .A(n42), .B(n60), .Z(n1166) );
  AO7SVTX2 U1721 ( .A(n1794), .B(n136), .C(n1793), .Z(n1795) );
  F_ND2SVTX1 U1722 ( .A(n1840), .B(n110), .Z(n1773) );
  AO6SVTX2 U1723 ( .A(n1842), .B(n110), .C(n1841), .Z(n1843) );
  ENSVTX0H U1724 ( .A(n1500), .B(n1499), .Z(n1512) );
  IVSVTX4 U1725 ( .A(n1827), .Z(n907) );
  IVSVTX2 U1726 ( .A(n1631), .Z(n745) );
  IVSVTX2 U1727 ( .A(n980), .Z(n764) );
  IVSVTX4 U1728 ( .A(n763), .Z(n1078) );
  AN2SVTX4 U1729 ( .A(n1041), .B(n1040), .Z(n805) );
  IVSVTX2 U1730 ( .A(n1034), .Z(n1035) );
  IVSVTX2 U1731 ( .A(n1228), .Z(n1220) );
  NR2SVTX2 U1732 ( .A(n1338), .B(n1282), .Z(n1281) );
  AO6SVTX2 U1733 ( .A(n69), .B(n499), .C(n1071), .Z(n1077) );
  NR2SVTX2 U1734 ( .A(n218), .B(n896), .Z(n1527) );
  AO7SVTX1 U1735 ( .A(n1690), .B(n1985), .C(n1689), .Z(n1691) );
  NR2SVTX2 U1736 ( .A(n1546), .B(n1906), .Z(n1549) );
  NR2SVTX0H U1737 ( .A(n2004), .B(n80), .Z(n2009) );
  NR2SVTX2 U1738 ( .A(n1858), .B(n1989), .Z(n1991) );
  AO7SVTX2 U1739 ( .A(n1878), .B(n1877), .C(n1876), .Z(n1879) );
  AO7NSVTX6 U1740 ( .A(n1902), .B(n1766), .C(n778), .Z(n780) );
  AO7SVTX2 U1741 ( .A(n939), .B(n895), .C(n896), .Z(n941) );
  F_ND2SVTX0H U1742 ( .A(n2017), .B(n2019), .Z(n1942) );
  ND2SVTX4 U1743 ( .A(n816), .B(n898), .Z(n2017) );
  ND2SVTX4 U1744 ( .A(m1[12]), .B(n889), .Z(n1506) );
  AO7SVTX4 U1745 ( .A(n738), .B(n1105), .C(n1519), .Z(n1092) );
  IVSVTX2 U1746 ( .A(n1038), .Z(n1042) );
  NR2SVTX2 U1747 ( .A(m1[23]), .B(n1053), .Z(n1056) );
  ND2SVTX2 U1748 ( .A(m1[23]), .B(n1025), .Z(n839) );
  ENSVTX4 U1749 ( .A(m1[23]), .B(n928), .Z(n972) );
  ND2SVTX2 U1750 ( .A(m1[8]), .B(n906), .Z(n1882) );
  ND2SVTX2 U1751 ( .A(n738), .B(n1792), .Z(n1703) );
  ND2SVTX2 U1752 ( .A(n954), .B(n354), .Z(n1270) );
  ND2SVTX2 U1753 ( .A(n928), .B(n354), .Z(n1218) );
  ND2SVTX2 U1754 ( .A(n759), .B(n938), .Z(n1719) );
  ND2SVTX4 U1755 ( .A(n62), .B(n1413), .Z(n1906) );
  ND2SVTX4 U1756 ( .A(n1188), .B(n1601), .Z(n1300) );
  ND2SVTX4 U1757 ( .A(n1358), .B(n1759), .Z(n1261) );
  ND2SVTX4 U1758 ( .A(n1519), .B(n1106), .Z(n2032) );
  ND2SVTX2 U1759 ( .A(n1543), .B(n1544), .Z(n1548) );
  OR2BSVTX6 U1760 ( .A(n889), .B(m1[17]), .Z(n1663) );
  ND2SVTX2 U1761 ( .A(n85), .B(n953), .Z(n1347) );
  OR2SVTX4 U1762 ( .A(n759), .B(n938), .Z(n776) );
  F_ND2SVTX0H U1763 ( .A(n1719), .B(n776), .Z(n1720) );
  ND2SVTX4 U1764 ( .A(n1475), .B(n776), .Z(n1580) );
  IVSVTX4 U1765 ( .A(n978), .Z(n979) );
  ND2SVTX2 U1766 ( .A(n758), .B(n1792), .Z(n1786) );
  ND2ASVTX8 U1767 ( .A(n1062), .B(n774), .Z(n1041) );
  ND2SVTX4 U1768 ( .A(n1192), .B(n1194), .Z(n956) );
  AO7SVTX4 U1769 ( .A(n895), .B(n1117), .C(n1927), .Z(n1521) );
  EOSVTX8 U1770 ( .A(n1253), .B(n1252), .Z(n769) );
  ND2SVTX2 U1771 ( .A(n1493), .B(n1494), .Z(n770) );
  NR2SVTX2 U1772 ( .A(n738), .B(n1123), .Z(n1694) );
  IVSVTX2 U1773 ( .A(n972), .Z(n973) );
  ND2SVTX2 U1774 ( .A(m1[25]), .B(n1068), .Z(n1022) );
  ND2SVTX2 U1775 ( .A(n1345), .B(m1[20]), .Z(n1331) );
  IVSVTX2 U1776 ( .A(n1555), .Z(n1030) );
  ND2SVTX2 U1777 ( .A(n171), .B(n85), .Z(n1631) );
  ND2SVTX4 U1778 ( .A(n1096), .B(n1095), .Z(n1682) );
  AO8SVTX2 U1779 ( .A(n1842), .B(n1498), .C(n172), .D(n1497), .Z(n1499) );
  ND2SVTX2 U1780 ( .A(n1663), .B(n1664), .Z(n1321) );
  AO8SVTX2 U1781 ( .A(n1842), .B(n1591), .C(n1451), .D(n1590), .Z(n1592) );
  B_ND2SVTX2 U1782 ( .A(n738), .B(n1105), .Z(n1093) );
  AO5SVTX2 U1783 ( .A(n1792), .B(n759), .C(m1[12]), .Z(n1135) );
  F_ENSVTX2 U1784 ( .A(n1629), .B(n1628), .Z(n1657) );
  AO8SVTX2 U1785 ( .A(n1842), .B(n187), .C(n1451), .D(n1626), .Z(n1628) );
  OR2SVTX4 U1786 ( .A(n56), .B(n55), .Z(n781) );
  NR2ASVTX2 U1787 ( .A(n672), .B(n355), .Z(n1051) );
  IVSVTX8 U1788 ( .A(m1[5]), .Z(n817) );
  F_ENSVTX2 U1789 ( .A(n1593), .B(n1592), .Z(n1611) );
  BFSVTX12 U1790 ( .A(n1485), .Z(n1670) );
  NR2SVTX2 U1791 ( .A(m1[23]), .B(n515), .Z(n1038) );
  ND2SVTX2 U1792 ( .A(n1569), .B(n1165), .Z(n1572) );
  ND2SVTX2 U1793 ( .A(m1[8]), .B(n758), .Z(n1861) );
  ND2SVTX4 U1794 ( .A(n1169), .B(n994), .Z(n1047) );
  AO5NSVTX4 U1795 ( .A(n1519), .B(n816), .C(n1116), .Z(n792) );
  AN2SVTX4 U1796 ( .A(m1[24]), .B(n1068), .Z(n1075) );
  IVSVTX8 U1797 ( .A(n1904), .Z(n1908) );
  ND2SVTX4 U1798 ( .A(n1854), .B(n1853), .Z(n1857) );
  AN2SVTX0H U1799 ( .A(m1[23]), .B(n666), .Z(n784) );
  OR2SVTX1 U1800 ( .A(n1038), .B(n999), .Z(n787) );
  F_AN2SVTX2 U1801 ( .A(n872), .B(n1157), .Z(n797) );
  BFSVTX2 U1802 ( .A(m1[26]), .Z(n968) );
  F_EOSVTX2 U1803 ( .A(n1290), .B(n1289), .Z(n800) );
  AN2SVTX0H U1804 ( .A(n712), .B(n1304), .Z(n804) );
  IVSVTX4 U1805 ( .A(n1086), .Z(n872) );
  OR2SVTX4 U1806 ( .A(n1755), .B(n921), .Z(n808) );
  IVSVTX2 U1807 ( .A(n1400), .Z(n943) );
  IVSVTX2 U1808 ( .A(n945), .Z(n1709) );
  F_ND2ASVTX2 U1809 ( .A(n944), .B(n1116), .Z(n945) );
  ND2ASVTX8 U1810 ( .A(n682), .B(n1975), .Z(n1399) );
  NR2ASVTX6 U1811 ( .A(n293), .B(n928), .Z(n1285) );
  ND2SVTX4 U1812 ( .A(m1[24]), .B(n196), .Z(n978) );
  ND2ASVTX8 U1813 ( .A(n889), .B(n708), .Z(n1642) );
  NR2SVTX4 U1814 ( .A(m1[10]), .B(n1102), .Z(n1964) );
  NR2SVTX4 U1815 ( .A(n1964), .B(n1972), .Z(n837) );
  NR2SVTX2 U1816 ( .A(n2044), .B(n1395), .Z(n1704) );
  ND2SVTX4 U1817 ( .A(n837), .B(n1704), .Z(n1446) );
  IVSVTX4 U1818 ( .A(n1396), .Z(n838) );
  ND2SVTX4 U1819 ( .A(n1519), .B(n1105), .Z(n2045) );
  AO7SVTX4 U1820 ( .A(n2045), .B(n1395), .C(n1393), .Z(n1969) );
  ND2SVTX4 U1821 ( .A(n1102), .B(n462), .Z(n1966) );
  IVSVTX4 U1822 ( .A(n844), .Z(n846) );
  IVSVTX4 U1823 ( .A(n1801), .Z(n858) );
  NR2SVTX6 U1824 ( .A(n273), .B(n734), .Z(n2015) );
  NR2SVTX4 U1825 ( .A(n2015), .B(n1941), .Z(n1372) );
  ND2SVTX6 U1826 ( .A(n866), .B(n865), .Z(n1696) );
  ND2SVTX4 U1827 ( .A(n1481), .B(n1480), .Z(n1614) );
  NR2SVTX4 U1828 ( .A(n928), .B(n1000), .Z(n1156) );
  NR2SVTX4 U1829 ( .A(n1068), .B(n515), .Z(n1083) );
  ND2SVTX4 U1830 ( .A(n76), .B(n917), .Z(n1206) );
  ND2SVTX2 U1831 ( .A(n605), .B(n515), .Z(n1085) );
  ND2SVTX8 U1832 ( .A(n1188), .B(n915), .Z(n1357) );
  IVSVTX4 U1833 ( .A(n1041), .Z(n1039) );
  IVSVTX4 U1834 ( .A(n891), .Z(n893) );
  ND2SVTX4 U1835 ( .A(n1519), .B(n896), .Z(n2052) );
  NR2ASVTX8 U1836 ( .A(n715), .B(n273), .Z(n2049) );
  NR2SVTX6 U1837 ( .A(n2056), .B(n2049), .Z(n899) );
  ND2SVTX4 U1838 ( .A(n2052), .B(n899), .Z(n901) );
  IVSVTX2 U1839 ( .A(n1527), .Z(n897) );
  ND2ASVTX6 U1840 ( .A(n715), .B(n273), .Z(n2051) );
  NR2SVTX4 U1841 ( .A(n758), .B(n1792), .Z(n902) );
  ND2SVTX8 U1842 ( .A(n794), .B(n910), .Z(n1320) );
  ND2SVTX4 U1843 ( .A(n923), .B(n922), .Z(n976) );
  ND2SVTX2 U1844 ( .A(n976), .B(n975), .Z(n1419) );
  NR2ASVTX8 U1845 ( .A(n927), .B(n926), .Z(n1279) );
  FAS1SVTX4 U1846 ( .A(n666), .B(n347), .CI(n1068), .CO(n923), .Z(n929) );
  ND2SVTX4 U1847 ( .A(n930), .B(n929), .Z(n1189) );
  ND2SVTX4 U1848 ( .A(n954), .B(n99), .Z(n994) );
  NR2SVTX2 U1849 ( .A(n716), .B(n1934), .Z(n1928) );
  NR2SVTX2 U1850 ( .A(n738), .B(n716), .Z(n1400) );
  ND2SVTX4 U1851 ( .A(n1775), .B(n856), .Z(n1958) );
  ND2SVTX2 U1852 ( .A(n917), .B(n928), .Z(n1193) );
  ND2SVTX4 U1853 ( .A(n1168), .B(n957), .Z(n959) );
  IVSVTX2 U1854 ( .A(n959), .Z(n955) );
  F_ND2ASVTX2 U1855 ( .A(m1[16]), .B(n708), .Z(n1759) );
  AO7ABSVTX4 U1856 ( .A(n46), .B(n959), .C(n958), .Z(n963) );
  ND2SVTX4 U1857 ( .A(n974), .B(n973), .Z(n1555) );
  B_ND2SVTX2 U1858 ( .A(n1180), .B(n61), .Z(n984) );
  NR2ASVTX6 U1859 ( .A(n178), .B(n1047), .Z(n996) );
  ND2SVTX4 U1860 ( .A(n996), .B(n1173), .Z(n1011) );
  NR2ASVTX6 U1861 ( .A(n1016), .B(n1015), .Z(n1018) );
  IVSVTX2 U1862 ( .A(n1022), .Z(n1082) );
  ND2SVTX4 U1863 ( .A(n1024), .B(n1023), .Z(n1029) );
  NR2ASVTX2 U1864 ( .A(m1[23]), .B(n1601), .Z(n1032) );
  ND2SVTX4 U1865 ( .A(n1554), .B(n1030), .Z(n1545) );
  ND2SVTX4 U1866 ( .A(n1052), .B(n1051), .Z(n1058) );
  IVSVTX0H U1867 ( .A(n1083), .Z(n1084) );
  NR2SVTX2 U1868 ( .A(n1156), .B(n649), .Z(n1087) );
  NR2SVTX4 U1869 ( .A(n777), .B(n1090), .Z(n1338) );
  NR2SVTX4 U1870 ( .A(n1279), .B(n1338), .Z(n1413) );
  FAS1SVTX4 U1871 ( .A(n682), .B(m1[8]), .CI(n1094), .CO(n1096), .Z(n1383) );
  IVSVTX4 U1872 ( .A(n1681), .Z(n1097) );
  IVSVTX4 U1873 ( .A(n1122), .Z(n1112) );
  ND2SVTX2 U1874 ( .A(n1110), .B(n1109), .Z(n2063) );
  AO7SVTX8 U1875 ( .A(n2062), .B(n2010), .C(n2063), .Z(n1390) );
  ND3SVTX8 U1876 ( .A(n1112), .B(n1390), .C(n1121), .Z(n1325) );
  ND2SVTX4 U1877 ( .A(n1114), .B(n1113), .Z(n2011) );
  FAS1SVTX4 U1878 ( .A(n222), .B(n751), .CI(n244), .CO(n1133), .Z(n1493) );
  ND2SVTX2 U1879 ( .A(n889), .B(n244), .Z(n1129) );
  ND2SVTX6 U1880 ( .A(n1341), .B(n1340), .Z(n1146) );
  ND2SVTX8 U1881 ( .A(n1543), .B(n1544), .Z(n1904) );
  IVSVTX0H U1882 ( .A(n1156), .Z(n1157) );
  IVSVTX0H U1883 ( .A(n788), .Z(n1183) );
  IVSVTX2 U1884 ( .A(n1185), .Z(n1205) );
  ND2SVTX4 U1885 ( .A(n1422), .B(n1420), .Z(n1187) );
  NR2SVTX6 U1886 ( .A(n1187), .B(n1423), .Z(n1211) );
  ND2SVTX2 U1887 ( .A(n1193), .B(n1192), .Z(n1196) );
  NR2ASVTX2 U1888 ( .A(n1196), .B(n1197), .Z(n1201) );
  IVSVTX2 U1889 ( .A(n1196), .Z(n1199) );
  NR2SVTX2 U1890 ( .A(n1217), .B(n1216), .Z(n1226) );
  IVSVTX0H U1891 ( .A(n919), .Z(n1223) );
  IVSVTX2 U1892 ( .A(n1221), .Z(n1222) );
  F_ND2ASVTX2 U1893 ( .A(n1223), .B(n1222), .Z(n1236) );
  IVSVTX2 U1894 ( .A(n1226), .Z(n1231) );
  NR3SVTX2 U1895 ( .A(n1231), .B(n1228), .C(n163), .Z(n1229) );
  ND3SVTX2 U1896 ( .A(n320), .B(n1229), .C(n1230), .Z(n1235) );
  IVSVTX2 U1897 ( .A(n1230), .Z(n1233) );
  NR2ASVTX1 U1898 ( .A(n1231), .B(n163), .Z(n1232) );
  NR2SVTX4 U1899 ( .A(n1237), .B(n152), .Z(n1238) );
  NR2ASVTX6 U1900 ( .A(n706), .B(n1239), .Z(n1240) );
  ND3ABSVTX2 U1901 ( .A(n1258), .B(n1259), .C(n920), .Z(n1269) );
  IVSVTX0H U1902 ( .A(n1261), .Z(n1264) );
  IVSVTX0H U1903 ( .A(n1262), .Z(n1263) );
  IVSVTX4 U1904 ( .A(n1363), .Z(n1267) );
  IVSVTX4 U1905 ( .A(n756), .Z(n1275) );
  ND2ASVTX8 U1906 ( .A(n730), .B(n21), .Z(n1272) );
  IVSVTX4 U1907 ( .A(n1660), .Z(n1348) );
  NR2SVTX2 U1908 ( .A(n1272), .B(n1348), .Z(n1273) );
  NR2SVTX2 U1909 ( .A(n1285), .B(n1284), .Z(n1290) );
  NR2SVTX4 U1910 ( .A(n1306), .B(n1348), .Z(n1307) );
  ND2SVTX4 U1911 ( .A(n1316), .B(n1451), .Z(n1748) );
  IVSVTX4 U1912 ( .A(n1748), .Z(n1311) );
  IVSVTX4 U1913 ( .A(n452), .Z(n1309) );
  IVSVTX4 U1914 ( .A(n1277), .Z(n1364) );
  ND2SVTX2 U1915 ( .A(n1371), .B(n861), .Z(n1381) );
  NR2SVTX2 U1916 ( .A(n1373), .B(n2037), .Z(n1379) );
  AO7SVTX1 U1917 ( .A(n2037), .B(n1377), .C(n2039), .Z(n1378) );
  F_ND2ASVTX2 U1918 ( .A(n1387), .B(n1386), .Z(n2066) );
  ENSVTX0H U1919 ( .A(n1391), .B(n1856), .Z(n1392) );
  NR2SVTX2 U1920 ( .A(n1392), .B(n1902), .Z(n1410) );
  IVSVTX0H U1921 ( .A(n1393), .Z(n1394) );
  AO7SVTX1 U1922 ( .A(n2044), .B(n2046), .C(n2045), .Z(n1397) );
  ENSVTX0H U1923 ( .A(n1398), .B(n1397), .Z(n1408) );
  NR2ASVTX1 U1924 ( .A(n1399), .B(n1709), .Z(n1405) );
  IVSVTX0H U1925 ( .A(n2032), .Z(n1403) );
  AO6SVTX1 U1926 ( .A(n943), .B(n2033), .C(n1403), .Z(n1404) );
  ENSVTX0H U1927 ( .A(n1405), .B(n1404), .Z(n1406) );
  ND2SVTX4 U1928 ( .A(n815), .B(n1412), .Z(m2[4]) );
  BFSVTX1 U1929 ( .A(n1436), .Z(n1581) );
  AO6SVTX1 U1930 ( .A(n1435), .B(n1437), .C(n214), .Z(n1438) );
  AO7SVTX6 U1931 ( .A(n137), .B(n2046), .C(n1445), .Z(n1870) );
  AO7SVTX1 U1932 ( .A(n1651), .B(n216), .C(n1506), .Z(n1447) );
  F_ENSVTX2 U1933 ( .A(n1455), .B(n1454), .Z(n1456) );
  IVSVTX0H U1934 ( .A(n1457), .Z(n1459) );
  AO7SVTX2 U1935 ( .A(n1463), .B(n1461), .C(n1462), .Z(n1464) );
  AO8SVTX2 U1936 ( .A(n1603), .B(n139), .C(n1873), .D(n1464), .Z(n1465) );
  AO7ABSVTX4 U1937 ( .A(n1485), .B(n1473), .C(n1472), .Z(m2[12]) );
  AO6SVTX1 U1938 ( .A(n1435), .B(n776), .C(n1476), .Z(n1477) );
  EOSVTX0H U1939 ( .A(n1478), .B(n1477), .Z(n1489) );
  AO6SVTX1 U1940 ( .A(n219), .B(n1481), .C(n1482), .Z(n1483) );
  EOSVTX2 U1941 ( .A(n1484), .B(n1483), .Z(n1486) );
  BFSVTX6 U1942 ( .A(n1495), .Z(n1728) );
  AO7SVTX1 U1943 ( .A(n1727), .B(n1496), .C(n770), .Z(n1497) );
  ENSVTX0H U1944 ( .A(n1503), .B(n1502), .Z(n1504) );
  ENSVTX0H U1945 ( .A(n1508), .B(n1507), .Z(n1509) );
  ENSVTX0H U1946 ( .A(n1518), .B(n1927), .Z(n1514) );
  IVSVTX0H U1947 ( .A(n1931), .Z(n1515) );
  ENSVTX0H U1948 ( .A(n1933), .B(n1516), .Z(n1523) );
  AO7SVTX1 U1949 ( .A(n528), .B(n1518), .C(n1517), .Z(n1520) );
  ENSVTX0H U1950 ( .A(n1521), .B(n1520), .Z(n1522) );
  EOSVTX0H U1951 ( .A(n1527), .B(n1526), .Z(n1533) );
  ND2SVTX2 U1952 ( .A(n1528), .B(n1529), .Z(n1530) );
  EOSVTX0H U1953 ( .A(n1531), .B(n1530), .Z(n1532) );
  ND3SVTX4 U1954 ( .A(n1536), .B(n1535), .C(n1534), .Z(m2[0]) );
  ND2SVTX4 U1955 ( .A(n1555), .B(n1561), .Z(n1563) );
  NR3SVTX6 U1956 ( .A(n1560), .B(n1559), .C(n152), .Z(n1562) );
  ND3ABSVTX8 U1957 ( .A(n1919), .B(n1574), .C(n1573), .Z(n1924) );
  AO7SVTX1 U1958 ( .A(n1582), .B(n1581), .C(n419), .Z(n1583) );
  AO6SVTX2 U1959 ( .A(n1435), .B(n1584), .C(n1583), .Z(n1585) );
  F_EOSVTX2 U1960 ( .A(n1586), .B(n1585), .Z(n1622) );
  IVSVTX0H U1961 ( .A(n1588), .Z(n1589) );
  IVSVTX0H U1962 ( .A(n1643), .Z(n1595) );
  IVSVTX0H U1963 ( .A(n1646), .Z(n1594) );
  AO7SVTX1 U1964 ( .A(n1595), .B(n212), .C(n1594), .Z(n1596) );
  ENSVTX0H U1965 ( .A(n1599), .B(n1598), .Z(n1600) );
  NR2SVTX2 U1966 ( .A(n1600), .B(n1877), .Z(n1610) );
  NR3ABSVTX2 U1967 ( .A(n1603), .B(n66), .C(n1636), .Z(n1605) );
  AO7SVTX1 U1968 ( .A(n1461), .B(n739), .C(n27), .Z(n1604) );
  NR2SVTX2 U1969 ( .A(n1605), .B(n1604), .Z(n1606) );
  AO4SVTX1 U1970 ( .A(n44), .B(n675), .C(n1608), .D(n60), .Z(n1609) );
  ND2SVTX1 U1971 ( .A(n1613), .B(n444), .Z(n1619) );
  NR2SVTX2 U1972 ( .A(n1615), .B(n1614), .Z(n1617) );
  IVSVTX0H U1973 ( .A(n1623), .Z(n1624) );
  AO7SVTX1 U1974 ( .A(n749), .B(n27), .C(n138), .Z(n1633) );
  AO6ABSVTX2 U1975 ( .A(n1461), .B(n1635), .C(n1633), .Z(n1634) );
  IVSVTX0H U1976 ( .A(n1644), .Z(n1645) );
  AO6SVTX1 U1977 ( .A(n1646), .B(n17), .C(n1645), .Z(n1648) );
  ENSVTX0H U1978 ( .A(n1653), .B(n1652), .Z(n1654) );
  AO6SVTX1 U1979 ( .A(n219), .B(n1660), .C(n1659), .Z(n1661) );
  ND2ASVTX8 U1980 ( .A(n1671), .B(n813), .Z(m2[14]) );
  IVSVTX4 U1981 ( .A(n2080), .Z(n1679) );
  NR2ASVTX6 U1982 ( .A(n771), .B(n1677), .Z(n2077) );
  AO6CSVTX8 U1983 ( .A(n2076), .B(n1679), .C(n1678), .Z(n1898) );
  EOSVTX8 U1984 ( .A(n1680), .B(n1898), .Z(m2[17]) );
  ENSVTX0H U1985 ( .A(n1692), .B(n1691), .Z(n1693) );
  IVSVTX0H U1986 ( .A(n1694), .Z(n1695) );
  IVSVTX2 U1987 ( .A(n1696), .Z(n1954) );
  EOSVTX0H U1988 ( .A(n1697), .B(n1954), .Z(n1698) );
  NR2SVTX2 U1989 ( .A(n1967), .B(n737), .Z(n1707) );
  IVSVTX0H U1990 ( .A(n1704), .Z(n1971) );
  AO7SVTX1 U1991 ( .A(n1971), .B(n2046), .C(n1705), .Z(n1706) );
  ENSVTX0H U1992 ( .A(n1707), .B(n1706), .Z(n1715) );
  IVSVTX0H U1993 ( .A(n1710), .Z(n1711) );
  AO1CDSVTX2 U1994 ( .A(n2033), .B(n782), .C(n945), .D(n1711), .Z(n1960) );
  ENSVTX0H U1995 ( .A(n1712), .B(n1960), .Z(n1713) );
  ND2SVTX2 U1996 ( .A(n1481), .B(n1717), .Z(n1718) );
  ENSVTX0H U1997 ( .A(n1720), .B(n1435), .Z(n1745) );
  ND2SVTX2 U1998 ( .A(n1722), .B(n1721), .Z(n1726) );
  AO7SVTX1 U1999 ( .A(n1723), .B(n1814), .C(n1813), .Z(n1724) );
  AO8SVTX1 U2000 ( .A(n1816), .B(n1812), .C(n1870), .D(n1724), .Z(n1725) );
  ENSVTX0H U2001 ( .A(n1726), .B(n1725), .Z(n1743) );
  NR2ASVTX1 U2002 ( .A(n770), .B(n1727), .Z(n1731) );
  AO6SVTX2 U2003 ( .A(n1842), .B(n172), .C(n1728), .Z(n1730) );
  F_ENSVTX2 U2004 ( .A(n1731), .B(n1730), .Z(n1732) );
  AO7SVTX1 U2005 ( .A(n1819), .B(n1734), .C(n1125), .Z(n1736) );
  AO7SVTX6 U2006 ( .A(n921), .B(n810), .C(n1746), .Z(m2[10]) );
  NR2ASVTX1 U2007 ( .A(n1751), .B(n1750), .Z(n1752) );
  F_ENSVTX2 U2008 ( .A(n1761), .B(n353), .Z(n1762) );
  AO7SVTX1 U2009 ( .A(n158), .B(n1954), .C(n18), .Z(n1770) );
  ENSVTX0H U2010 ( .A(n1771), .B(n1770), .Z(n1772) );
  ENSVTX0H U2011 ( .A(n1780), .B(n1779), .Z(n1798) );
  NR2ASVTX1 U2012 ( .A(n1781), .B(n87), .Z(n1785) );
  AO6SVTX1 U2013 ( .A(n1873), .B(n1872), .C(n937), .Z(n1784) );
  ENSVTX0H U2014 ( .A(n1785), .B(n1784), .Z(n1796) );
  AO7SVTX2 U2015 ( .A(n1985), .B(n190), .C(n164), .Z(n1789) );
  ENSVTX0H U2016 ( .A(n1790), .B(n1789), .Z(n1791) );
  F_IVSVTX1 U2017 ( .A(n158), .Z(n1803) );
  AO6SVTX1 U2018 ( .A(n1805), .B(n409), .C(n1804), .Z(n1806) );
  AO7SVTX1 U2019 ( .A(n1954), .B(n1807), .C(n1806), .Z(n1808) );
  ENSVTX0H U2020 ( .A(n1809), .B(n1808), .Z(n1810) );
  AO6SVTX1 U2021 ( .A(n1870), .B(n1816), .C(n1815), .Z(n1817) );
  ENSVTX0H U2022 ( .A(n1818), .B(n1817), .Z(n1825) );
  NR2ASVTX1 U2023 ( .A(n1125), .B(n1734), .Z(n1822) );
  ENSVTX0H U2024 ( .A(n1822), .B(n1821), .Z(n1823) );
  ND2SVTX2 U2025 ( .A(n1828), .B(n1827), .Z(n1836) );
  IVSVTX0H U2026 ( .A(n164), .Z(n1832) );
  AO6SVTX1 U2027 ( .A(n1832), .B(n1831), .C(n1830), .Z(n1833) );
  ENSVTX0H U2028 ( .A(n1836), .B(n1835), .Z(n1846) );
  NR2SVTX2 U2029 ( .A(n1854), .B(n1853), .Z(n1989) );
  AO7SVTX2 U2030 ( .A(n1989), .B(n1990), .C(n1857), .Z(n1859) );
  IVSVTX0H U2031 ( .A(n1863), .Z(n1866) );
  AO7SVTX1 U2032 ( .A(n1866), .B(n1954), .C(n1865), .Z(n1867) );
  ENSVTX0H U2033 ( .A(n1868), .B(n1867), .Z(n1880) );
  NR2ASVTX1 U2034 ( .A(n217), .B(n3), .Z(n1871) );
  ENSVTX0H U2035 ( .A(n1871), .B(n1870), .Z(n1878) );
  ENSVTX0H U2036 ( .A(n1874), .B(n1873), .Z(n1875) );
  AO7SVTX1 U2037 ( .A(n1889), .B(n1985), .C(n1888), .Z(n1890) );
  ENSVTX0H U2038 ( .A(n1891), .B(n1890), .Z(n1892) );
  AO3SVTX4 U2039 ( .A(n1902), .B(n1895), .C(n1894), .D(n1893), .Z(m2[7]) );
  IVSVTX2 U2040 ( .A(n1897), .Z(n1899) );
  AO7SVTX6 U2041 ( .A(n1899), .B(n1898), .C(n723), .Z(n1900) );
  ENSVTX0H U2042 ( .A(n1999), .B(n1929), .Z(n1930) );
  AO7SVTX1 U2043 ( .A(n1933), .B(n1932), .C(n1931), .Z(n2007) );
  ENSVTX0H U2044 ( .A(n2007), .B(n1936), .Z(n1940) );
  ND2SVTX2 U2045 ( .A(n705), .B(n1385), .Z(n1937) );
  ENSVTX0H U2046 ( .A(n1938), .B(n1937), .Z(n1939) );
  ENSVTX0H U2047 ( .A(n1942), .B(n2040), .Z(n1943) );
  ENSVTX0H U2048 ( .A(n2058), .B(n1945), .Z(n1946) );
  ND2SVTX2 U2049 ( .A(n1953), .B(n1952), .Z(n1956) );
  ENSVTX0H U2050 ( .A(n1956), .B(n1955), .Z(n1981) );
  ENSVTX0H U2051 ( .A(n1963), .B(n1962), .Z(n1979) );
  IVSVTX0H U2052 ( .A(n1964), .Z(n1965) );
  IVSVTX0H U2053 ( .A(n737), .Z(n1968) );
  AO6SVTX1 U2054 ( .A(n1969), .B(n1968), .C(n1967), .Z(n1970) );
  AO21SVTX1 U2055 ( .A(n737), .B(n1971), .C(n2046), .D(n1970), .Z(n1973) );
  ENSVTX0H U2056 ( .A(n1974), .B(n1973), .Z(n1976) );
  AO2ABSVTX1 U2057 ( .C(n1976), .D(n37), .A(n1975), .B(n44), .Z(n1977) );
  AO7SVTX1 U2058 ( .A(n1986), .B(n1985), .C(n1984), .Z(n1987) );
  ENSVTX0H U2059 ( .A(n1988), .B(n1987), .Z(n1993) );
  ENSVTX0H U2060 ( .A(n1991), .B(n1990), .Z(n1992) );
  NR2SVTX2 U2061 ( .A(n1995), .B(n762), .Z(n2001) );
  IVSVTX0H U2062 ( .A(n1996), .Z(n1997) );
  AO6SVTX1 U2063 ( .A(n1999), .B(n1998), .C(n1997), .Z(n2000) );
  ENSVTX0H U2064 ( .A(n2001), .B(n2000), .Z(n2002) );
  IVSVTX0H U2065 ( .A(n2005), .Z(n2006) );
  AO6SVTX1 U2066 ( .A(n2007), .B(n88), .C(n2006), .Z(n2008) );
  ENSVTX0H U2067 ( .A(n2009), .B(n2008), .Z(n2014) );
  F_ND2ASVTX2 U2068 ( .A(n2064), .B(n2065), .Z(n2012) );
  ENSVTX0H U2069 ( .A(n2012), .B(n2066), .Z(n2013) );
  F_AO2SVTX1 U2070 ( .A(n36), .B(n2014), .C(n174), .D(n2013), .Z(n2030) );
  AO6SVTX1 U2071 ( .A(n2058), .B(n2052), .C(n2024), .Z(n2025) );
  EOSVTX0H U2072 ( .A(n2026), .B(n2025), .Z(n2027) );
  ENSVTX0H U2073 ( .A(n2034), .B(n2033), .Z(n2035) );
  ENSVTX0H U2074 ( .A(n2047), .B(n2046), .Z(n2048) );
  AO7SVTX1 U2075 ( .A(n2056), .B(n2055), .C(n2054), .Z(n2057) );
  AO6SVTX1 U2076 ( .A(n2059), .B(n2058), .C(n2057), .Z(n2060) );
  EOSVTX0H U2077 ( .A(n2061), .B(n2060), .Z(n2070) );
  AO6SVTX1 U2078 ( .A(n2066), .B(n2065), .C(n2064), .Z(n2067) );
  ENSVTX0H U2079 ( .A(n2068), .B(n2067), .Z(n2069) );
  IVSVTX2 U2080 ( .A(n2076), .Z(n2078) );
  NR2SVTX2 U2081 ( .A(n2078), .B(n2077), .Z(n2079) );
  ENSVTX4 U2082 ( .A(n2080), .B(n2079), .Z(m2[16]) );
endmodule


module remap_top ( num_i, rslt_o );
  input [31:0] num_i;
  output [31:0] rslt_o;
  wire   n167, n169, n170, n171, n172, n173, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n217, n218, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n230, n231, n232, n233, n234, n235, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n359, n360, n361, n362, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728;
  wire   [27:0] keyvalues_m1;

  remap re_map ( .m1({keyvalues_m1[27:26], n180, n470, keyvalues_m1[23:21], 
        n445, keyvalues_m1[19:0]}), .m2(rslt_o[26:0]) );
  BFSVTX0H U200 ( .A(n718), .Z(rslt_o[30]) );
  IVSVTX10 U201 ( .A(n335), .Z(n470) );
  IVSVTX2 U202 ( .A(n239), .Z(n238) );
  IVSVTX2 U203 ( .A(n560), .Z(n563) );
  IVSVTX8 U204 ( .A(n566), .Z(keyvalues_m1[1]) );
  AO7CSVTX6 U205 ( .A(n386), .B(n428), .C(n246), .Z(n338) );
  ND3SVTX4 U206 ( .A(n359), .B(n360), .C(n299), .Z(n441) );
  ND3SVTX4 U207 ( .A(n385), .B(n693), .C(n712), .Z(n461) );
  NR3SVTX6 U208 ( .A(rslt_o[29]), .B(rslt_o[28]), .C(n293), .Z(n535) );
  IVSVTX2 U209 ( .A(n636), .Z(n293) );
  IVSVTX2 U210 ( .A(n416), .Z(n186) );
  IVSVTX8 U211 ( .A(n466), .Z(rslt_o[27]) );
  IVSVTX6 U212 ( .A(n277), .Z(rslt_o[28]) );
  ND3SVTX6 U213 ( .A(n725), .B(n693), .C(n724), .Z(n666) );
  B_ND2SVTX2 U214 ( .A(n201), .B(n634), .Z(n426) );
  AO2SVTX4 U215 ( .A(n284), .B(n687), .C(n181), .D(n396), .Z(n638) );
  ND2ASVTX6 U216 ( .A(n305), .B(n573), .Z(n574) );
  IVSVTX2 U217 ( .A(n720), .Z(n554) );
  IVSVTX8 U218 ( .A(n246), .Z(n687) );
  ND2ASVTX4 U219 ( .A(n408), .B(n639), .Z(n713) );
  ND2SVTX4 U220 ( .A(n592), .B(n593), .Z(n385) );
  ND2SVTX2 U221 ( .A(n396), .B(n685), .Z(n541) );
  BFSVTX2 U222 ( .A(n364), .Z(n201) );
  CTBUFSVTX4 U223 ( .A(n414), .Z(n225) );
  AO7SVTX2 U224 ( .A(n561), .B(n345), .C(n600), .Z(n348) );
  CTIVSVTX2 U225 ( .A(n249), .Z(n452) );
  IVSVTX6 U226 ( .A(n709), .Z(n396) );
  IVSVTX4 U227 ( .A(n693), .Z(n417) );
  AN2SVTX6 U228 ( .A(n464), .B(n304), .Z(n416) );
  IVSVTX2 U229 ( .A(n695), .Z(n311) );
  AO2SVTX6 U230 ( .A(n383), .B(n685), .C(n259), .D(n187), .Z(n260) );
  AO2SVTX4 U231 ( .A(n594), .B(n585), .C(n453), .D(n677), .Z(n723) );
  AO7SVTX2 U232 ( .A(n401), .B(n611), .C(n624), .Z(n612) );
  NR2SVTX4 U233 ( .A(n283), .B(n589), .Z(n710) );
  IVSVTX6 U234 ( .A(n271), .Z(n272) );
  CTIVSVTX6 U235 ( .A(n383), .Z(n199) );
  IVSVTX2 U236 ( .A(n583), .Z(n248) );
  AO7SVTX1 U237 ( .A(n606), .B(n301), .C(n605), .Z(n607) );
  NR2ASVTX2 U238 ( .A(n610), .B(n228), .Z(n611) );
  NR2SVTX6 U239 ( .A(n691), .B(n279), .Z(n259) );
  IVSVTX2 U240 ( .A(n406), .Z(n705) );
  ND3SVTX4 U241 ( .A(n667), .B(n464), .C(n365), .Z(n695) );
  AO20SVTX4 U242 ( .A(n191), .B(n618), .C(n193), .D(rslt_o[31]), .Z(n621) );
  IVSVTX6 U243 ( .A(n228), .Z(n187) );
  IVSVTX8 U244 ( .A(n279), .Z(n364) );
  IVSVTX2 U245 ( .A(n691), .Z(n366) );
  CTIVSVTX4 U246 ( .A(n718), .Z(n345) );
  IVSVTX10 U247 ( .A(n274), .Z(n383) );
  NR2ASVTX4 U248 ( .A(num_i[13]), .B(n559), .Z(n352) );
  AO7SVTX4 U249 ( .A(n481), .B(rslt_o[31]), .C(n267), .Z(n266) );
  IVSVTX0H U250 ( .A(n526), .Z(n450) );
  AO7SVTX4 U251 ( .A(n663), .B(n436), .C(n552), .Z(n583) );
  AO7SVTX2 U252 ( .A(n302), .B(n301), .C(n645), .Z(n667) );
  AO2ABSVTX6 U253 ( .C(n617), .D(n292), .A(n295), .B(n703), .Z(n294) );
  IVSVTX0H U254 ( .A(num_i[10]), .Z(n167) );
  IVSVTX6 U255 ( .A(n559), .Z(n292) );
  BFSVTX6 U256 ( .A(n471), .Z(n220) );
  IVSVTX0H U257 ( .A(n487), .Z(n588) );
  CTIVSVTX8 U258 ( .A(n365), .Z(n277) );
  NR2ASVTX4 U259 ( .A(n577), .B(n655), .Z(n692) );
  OR2SVTX2 U260 ( .A(n646), .B(n575), .Z(n302) );
  IVSVTX2 U261 ( .A(n446), .Z(n586) );
  BFSVTX2 U262 ( .A(num_i[4]), .Z(n706) );
  NR2ASVTX1 U263 ( .A(n567), .B(n183), .Z(n439) );
  AO7SVTX2 U264 ( .A(n659), .B(n658), .C(n327), .Z(n660) );
  IVSVTX0H U265 ( .A(num_i[25]), .Z(n267) );
  F_AN2SVTX2 U266 ( .A(num_i[13]), .B(n467), .Z(n658) );
  IVSVTX4 U267 ( .A(n609), .Z(n257) );
  IVSVTX2 U268 ( .A(n654), .Z(n468) );
  BFSVTX8 U269 ( .A(n663), .Z(n184) );
  NR2ASVTX4 U270 ( .A(n625), .B(n703), .Z(n568) );
  AO2SVTX4 U271 ( .A(n188), .B(n321), .C(n182), .D(n480), .Z(n241) );
  BFSVTX10 U272 ( .A(n411), .Z(n327) );
  B_ND2SVTX2 U273 ( .A(n647), .B(n471), .Z(n170) );
  NR2SVTX4 U274 ( .A(n258), .B(n288), .Z(n244) );
  F_ND2SVTX1 U275 ( .A(n657), .B(n309), .Z(n310) );
  NR2ASVTX4 U276 ( .A(n610), .B(n467), .Z(n579) );
  AN2SVTX1 U277 ( .A(num_i[13]), .B(n285), .Z(n480) );
  NR2ASVTX2 U278 ( .A(num_i[9]), .B(n703), .Z(n435) );
  BFSVTX2 U279 ( .A(num_i[6]), .Z(n567) );
  IVSVTX6 U280 ( .A(n522), .Z(n188) );
  NR3ABSVTX6 U281 ( .A(n525), .B(n412), .C(n326), .Z(n502) );
  BFSVTX2 U282 ( .A(num_i[7]), .Z(n610) );
  NR2SVTX4 U283 ( .A(n190), .B(n497), .Z(n258) );
  ND3SVTX4 U284 ( .A(n465), .B(n524), .C(n399), .Z(n357) );
  IVSVTX2 U285 ( .A(n538), .Z(n524) );
  F_ND2SVTX1 U286 ( .A(n646), .B(n514), .Z(n500) );
  AO7SVTX6 U287 ( .A(n603), .B(n484), .C(n189), .Z(n395) );
  IVSVTX2 U288 ( .A(num_i[3]), .Z(n728) );
  IVSVTX6 U289 ( .A(n413), .Z(n412) );
  IVSVTX2 U290 ( .A(n525), .Z(n505) );
  IVSVTX1 U291 ( .A(n520), .Z(n394) );
  IVSVTX4 U292 ( .A(n399), .Z(n508) );
  NR2SVTX2 U293 ( .A(n516), .B(n250), .Z(n391) );
  NR2SVTX6 U294 ( .A(n528), .B(n319), .Z(n375) );
  BFSVTX2 U295 ( .A(num_i[19]), .Z(n603) );
  CTBUFSVTX4 U296 ( .A(n331), .Z(n319) );
  IVSVTX4 U297 ( .A(n232), .Z(n525) );
  IVSVTX2 U298 ( .A(num_i[24]), .Z(n519) );
  IVSVTX2 U299 ( .A(num_i[14]), .Z(n285) );
  ND2SVTX2 U300 ( .A(n517), .B(n295), .Z(n250) );
  NR2SVTX2 U301 ( .A(num_i[7]), .B(num_i[6]), .Z(n514) );
  ND3SVTX4 U302 ( .A(num_i[19]), .B(n406), .C(n332), .Z(n173) );
  NR2SVTX2 U303 ( .A(num_i[11]), .B(num_i[10]), .Z(n373) );
  IVSVTX4 U304 ( .A(num_i[30]), .Z(n194) );
  BFSVTX4 U305 ( .A(num_i[26]), .Z(n529) );
  ND3SVTX4 U306 ( .A(num_i[15]), .B(n544), .C(n492), .Z(n489) );
  ND2SVTX6 U307 ( .A(n491), .B(n616), .Z(n490) );
  NR2SVTX4 U308 ( .A(num_i[21]), .B(num_i[20]), .Z(n387) );
  BFSVTX4 U309 ( .A(num_i[27]), .Z(n604) );
  IVSVTX4 U310 ( .A(num_i[31]), .Z(n456) );
  NR2SVTX2 U311 ( .A(num_i[5]), .B(num_i[4]), .Z(n513) );
  IVSVTX4 U312 ( .A(num_i[26]), .Z(n492) );
  CTIVSVTX4 U313 ( .A(n485), .Z(n486) );
  NR2SVTX4 U314 ( .A(num_i[22]), .B(num_i[23]), .Z(n231) );
  BFSVTX6 U315 ( .A(num_i[30]), .Z(n330) );
  ND4SVTX6 U316 ( .A(n359), .B(n360), .C(n693), .D(n299), .Z(n255) );
  ND2SVTX4 U317 ( .A(n249), .B(n397), .Z(n213) );
  AO7ABSVTX4 U318 ( .A(n651), .B(n354), .C(n650), .Z(n702) );
  NR3SVTX6 U319 ( .A(n693), .B(n312), .C(n311), .Z(n313) );
  IVSVTX4 U320 ( .A(n210), .Z(n397) );
  AO6SVTX8 U321 ( .A(n459), .B(n461), .C(n223), .Z(n460) );
  AO6SVTX6 U322 ( .A(n649), .B(n327), .C(n648), .Z(n662) );
  ND2SVTX2 U323 ( .A(n633), .B(n347), .Z(n329) );
  ND2SVTX4 U324 ( .A(n684), .B(n347), .Z(n337) );
  ND3SVTX8 U325 ( .A(n221), .B(n533), .C(n245), .Z(n340) );
  AO7CSVTX8 U326 ( .A(n535), .B(n340), .C(n466), .Z(n339) );
  IVSVTX6 U327 ( .A(n402), .Z(n172) );
  AO4SVTX6 U328 ( .A(n167), .B(n559), .C(n558), .D(n218), .Z(n639) );
  ND2SVTX4 U329 ( .A(n347), .B(n181), .Z(n215) );
  MUX21NSVTX8 U330 ( .A(n723), .B(n722), .S(n417), .Z(keyvalues_m1[3]) );
  ND2SVTX4 U331 ( .A(n652), .B(n656), .Z(n661) );
  ND2SVTX8 U332 ( .A(n636), .B(n383), .Z(n270) );
  ND2ASVTX8 U333 ( .A(n333), .B(n273), .Z(n670) );
  IVSVTX12 U334 ( .A(n257), .Z(n228) );
  AO4SVTX6 U335 ( .A(n228), .B(n692), .C(n464), .D(n691), .Z(n308) );
  ND2SVTX6 U336 ( .A(n693), .B(n382), .Z(n209) );
  IVSVTX8 U337 ( .A(n609), .Z(n464) );
  ND2ASVTX8 U338 ( .A(n609), .B(n306), .Z(n589) );
  NR3SVTX8 U339 ( .A(n463), .B(n598), .C(n184), .Z(n704) );
  IVSVTX4 U340 ( .A(n249), .Z(n169) );
  AO7ASVTX8 U341 ( .A(n169), .B(n717), .C(n680), .Z(keyvalues_m1[6]) );
  IVSVTX4 U342 ( .A(n170), .Z(n648) );
  ND2SVTX4 U343 ( .A(n228), .B(n367), .Z(n265) );
  OR3SVTX4 U344 ( .A(num_i[10]), .B(n481), .C(n497), .Z(n177) );
  BFSVTX12 U345 ( .A(n467), .Z(n301) );
  ND2ASVTX8 U346 ( .A(n413), .B(n399), .Z(n409) );
  AO3SVTX8 U347 ( .A(n522), .B(n390), .C(n171), .D(n626), .Z(n532) );
  ND3SVTX8 U348 ( .A(n399), .B(n412), .C(n518), .Z(n171) );
  IVSVTX12 U349 ( .A(n304), .Z(n305) );
  NR2SVTX6 U350 ( .A(num_i[18]), .B(num_i[19]), .Z(n483) );
  ND2SVTX6 U351 ( .A(n309), .B(n540), .Z(n507) );
  ND2SVTX4 U352 ( .A(n226), .B(n184), .Z(n590) );
  ND2SVTX4 U353 ( .A(n201), .B(n427), .Z(n615) );
  ND3SVTX6 U354 ( .A(n540), .B(n447), .C(n218), .Z(n230) );
  NR3SVTX8 U355 ( .A(n693), .B(n172), .C(n669), .Z(n424) );
  IVSVTX4 U356 ( .A(n173), .Z(n518) );
  AO7ABSVTX6 U357 ( .A(n367), .B(n690), .C(n307), .Z(n382) );
  IVSVTX12 U358 ( .A(n346), .Z(n347) );
  ND2SVTX4 U359 ( .A(n248), .B(n354), .Z(n298) );
  IVSVTX6 U360 ( .A(n211), .Z(n462) );
  AO4SVTX8 U361 ( .A(n277), .B(n281), .C(n278), .D(n279), .Z(n210) );
  ND2SVTX4 U362 ( .A(n657), .B(n471), .Z(n551) );
  F_ND2SVTX0H U363 ( .A(n705), .B(n601), .Z(n405) );
  ND2SVTX4 U364 ( .A(n396), .B(n635), .Z(n359) );
  ND2SVTX2 U365 ( .A(n185), .B(n193), .Z(n377) );
  IVSVTX2 U366 ( .A(n683), .Z(n328) );
  IVSVTX6 U367 ( .A(n506), .Z(n575) );
  OR2SVTX4 U368 ( .A(n718), .B(n619), .Z(n178) );
  AO7ABSVTX4 U369 ( .A(n220), .B(num_i[9]), .C(n660), .Z(n690) );
  AN2SVTX4 U370 ( .A(n687), .B(n681), .Z(n179) );
  MUX21NSVTX8 U371 ( .A(n689), .B(n688), .S(n687), .Z(n180) );
  MUX21SVTX8 U372 ( .A(n639), .B(n640), .S(n679), .Z(n181) );
  IVSVTX6 U373 ( .A(n212), .Z(n443) );
  AO2SVTX6 U374 ( .A(n347), .B(n636), .C(n415), .D(n434), .Z(n361) );
  CTBUFSVTX8 U375 ( .A(num_i[16]), .Z(n487) );
  AO2SVTX4 U376 ( .A(n602), .B(n464), .C(n601), .D(n220), .Z(n614) );
  IVSVTX12 U377 ( .A(n203), .Z(keyvalues_m1[17]) );
  IVSVTX12 U378 ( .A(n182), .Z(n183) );
  IVSVTX8 U379 ( .A(n208), .Z(n433) );
  ND4SVTX8 U380 ( .A(n596), .B(n394), .C(n419), .D(n399), .Z(n393) );
  IVSVTX10 U381 ( .A(n303), .Z(n419) );
  IVSVTX6 U382 ( .A(n400), .Z(n243) );
  IVSVTX8 U383 ( .A(n318), .Z(n182) );
  NR3SVTX4 U384 ( .A(n406), .B(n728), .C(n417), .Z(keyvalues_m1[0]) );
  ND3SVTX4 U385 ( .A(n185), .B(n193), .C(n233), .Z(n232) );
  ND2SVTX6 U386 ( .A(n557), .B(n556), .Z(n672) );
  AO7ABSVTX4 U387 ( .A(n685), .B(n416), .C(n337), .Z(n698) );
  IVSVTX8 U388 ( .A(n246), .Z(n466) );
  AO7SVTX2 U389 ( .A(n598), .B(n623), .C(n597), .Z(n599) );
  IVSVTX6 U390 ( .A(n187), .Z(rslt_o[29]) );
  ND2SVTX4 U391 ( .A(n718), .B(n439), .Z(n420) );
  ND2SVTX4 U392 ( .A(n608), .B(n586), .Z(n263) );
  IVSVTX8 U393 ( .A(n507), .Z(n663) );
  ND2ASVTX4 U394 ( .A(n349), .B(n197), .Z(n436) );
  NR3ABSVTX4 U395 ( .A(n193), .B(n285), .C(n523), .Z(n291) );
  CTIVSVTX4 U396 ( .A(n657), .Z(n598) );
  IVSVTX2 U397 ( .A(n521), .Z(n224) );
  B_ND2SVTX2 U398 ( .A(num_i[1]), .B(n498), .Z(n501) );
  IVSVTX2 U399 ( .A(n456), .Z(n457) );
  CTIVSVTX2 U400 ( .A(num_i[2]), .Z(n498) );
  IVSVTX4 U401 ( .A(num_i[8]), .Z(n191) );
  IVSVTX4 U402 ( .A(n632), .Z(n235) );
  NR2ASVTX6 U403 ( .A(n711), .B(n698), .Z(n336) );
  ND2SVTX6 U404 ( .A(n205), .B(n615), .Z(n239) );
  ND2SVTX6 U405 ( .A(n666), .B(n432), .Z(keyvalues_m1[11]) );
  NR2SVTX4 U406 ( .A(n186), .B(n276), .Z(n560) );
  ND2ASVTX4 U407 ( .A(n277), .B(n634), .Z(n681) );
  IVSVTX2 U408 ( .A(n699), .Z(n686) );
  IVSVTX8 U409 ( .A(n199), .Z(n273) );
  ND2SVTX4 U410 ( .A(n635), .B(n264), .Z(n261) );
  ND2SVTX6 U411 ( .A(n546), .B(n547), .Z(n386) );
  ND2SVTX6 U412 ( .A(n407), .B(n635), .Z(n712) );
  ND2SVTX6 U413 ( .A(n403), .B(n317), .Z(n669) );
  ND3SVTX4 U414 ( .A(n614), .B(n613), .C(n612), .Z(n427) );
  CTIVSVTX2 U415 ( .A(n623), .Z(n629) );
  ND2SVTX6 U416 ( .A(n420), .B(n437), .Z(n438) );
  IVSVTX2 U417 ( .A(n713), .Z(n715) );
  ND2SVTX6 U418 ( .A(n464), .B(n365), .Z(n709) );
  ND2SVTX6 U419 ( .A(n263), .B(n543), .Z(n635) );
  ND3ABSVTX8 U420 ( .A(n351), .B(n352), .C(n350), .Z(n685) );
  NR2ASVTX4 U421 ( .A(n596), .B(n718), .Z(n344) );
  NR2ASVTX4 U422 ( .A(num_i[11]), .B(n464), .Z(n401) );
  F_IVSVTX1 U423 ( .A(n633), .Z(n534) );
  B_ND2SVTX2 U424 ( .A(n627), .B(n626), .Z(n628) );
  ND2ASVTX4 U425 ( .A(n349), .B(n624), .Z(n561) );
  B_ND2SVTX2 U426 ( .A(n625), .B(n624), .Z(n627) );
  ND2SVTX4 U427 ( .A(n392), .B(n391), .Z(n390) );
  IVSVTX2 U428 ( .A(n290), .Z(n289) );
  AO6SVTX4 U429 ( .A(n515), .B(n514), .C(n377), .Z(n392) );
  B_ND2SVTX2 U430 ( .A(n706), .B(n705), .Z(n707) );
  NR3ABSVTX6 U431 ( .A(n519), .B(n520), .C(n224), .Z(n473) );
  IVSVTX6 U432 ( .A(n558), .Z(n455) );
  ND3SVTX4 U433 ( .A(n646), .B(n584), .C(n422), .Z(n421) );
  CTIVSVTX2 U434 ( .A(n610), .Z(n349) );
  NR2SVTX6 U435 ( .A(num_i[23]), .B(num_i[22]), .Z(n388) );
  NR2SVTX4 U436 ( .A(num_i[15]), .B(num_i[14]), .Z(n233) );
  IVSVTX4 U437 ( .A(num_i[10]), .Z(n192) );
  IVSVTX4 U438 ( .A(num_i[6]), .Z(n584) );
  IVSVTX4 U439 ( .A(num_i[18]), .Z(n558) );
  BFSVTX4 U440 ( .A(num_i[5]), .Z(n657) );
  IVSVTX8 U441 ( .A(num_i[9]), .Z(n481) );
  IVSVTX4 U442 ( .A(num_i[12]), .Z(n193) );
  IVSVTX6 U443 ( .A(num_i[13]), .Z(n185) );
  NR2SVTX4 U444 ( .A(n682), .B(n683), .Z(n689) );
  IVSVTX6 U445 ( .A(n671), .Z(n673) );
  ND2SVTX6 U446 ( .A(n261), .B(n260), .Z(n284) );
  NR2SVTX6 U447 ( .A(n669), .B(n315), .Z(n314) );
  IVSVTX4 U448 ( .A(n341), .Z(n245) );
  IVSVTX4 U449 ( .A(n549), .Z(n719) );
  AO6SVTX2 U450 ( .A(n629), .B(num_i[6]), .C(n628), .Z(n630) );
  IVSVTX4 U451 ( .A(n265), .Z(n264) );
  IVSVTX4 U452 ( .A(n333), .Z(n714) );
  NR2SVTX2 U453 ( .A(n344), .B(n595), .Z(n597) );
  IVSVTX4 U454 ( .A(n653), .Z(n278) );
  IVSVTX8 U455 ( .A(n300), .Z(n365) );
  ND3SVTX4 U456 ( .A(n652), .B(n282), .C(n468), .Z(n281) );
  IVSVTX4 U457 ( .A(n531), .Z(n251) );
  IVSVTX10 U458 ( .A(n408), .Z(n679) );
  AO7SVTX4 U459 ( .A(n655), .B(n654), .C(n327), .Z(n656) );
  IVSVTX2 U460 ( .A(n555), .Z(n384) );
  IVSVTX2 U461 ( .A(n537), .Z(n351) );
  AO6SVTX4 U462 ( .A(n463), .B(n455), .C(n529), .Z(n530) );
  IVSVTX4 U463 ( .A(n532), .Z(n252) );
  ND2SVTX4 U464 ( .A(n327), .B(n655), .Z(n282) );
  IVSVTX2 U465 ( .A(n202), .Z(n619) );
  IVSVTX2 U466 ( .A(n310), .Z(n659) );
  IVSVTX6 U467 ( .A(n411), .Z(n356) );
  NR4ABCSVTX6 U468 ( .A(n412), .B(n525), .C(n610), .D(n326), .Z(n321) );
  AO7SVTX6 U469 ( .A(n395), .B(n409), .C(n393), .Z(n400) );
  ND4ASVTX4 U470 ( .A(n538), .B(n525), .C(n378), .D(n379), .Z(n376) );
  ND4ABSVTX4 U471 ( .A(num_i[9]), .B(num_i[8]), .C(n423), .D(n421), .Z(n504)
         );
  NR2SVTX4 U472 ( .A(n325), .B(n324), .Z(n320) );
  ND2SVTX4 U473 ( .A(n494), .B(n495), .Z(n290) );
  IVSVTX8 U474 ( .A(n331), .Z(n189) );
  ND2SVTX6 U475 ( .A(n483), .B(n482), .Z(n538) );
  B_ND2SVTX2 U476 ( .A(num_i[5]), .B(n584), .Z(n499) );
  BFSVTX2 U477 ( .A(num_i[8]), .Z(n647) );
  BFSVTX2 U478 ( .A(num_i[12]), .Z(n617) );
  BFSVTX2 U479 ( .A(num_i[3]), .Z(n576) );
  NR2SVTX4 U480 ( .A(num_i[11]), .B(num_i[10]), .Z(n423) );
  NR2SVTX4 U481 ( .A(num_i[7]), .B(num_i[5]), .Z(n422) );
  IVSVTX6 U482 ( .A(num_i[4]), .Z(n646) );
  IVSVTX4 U483 ( .A(num_i[17]), .Z(n544) );
  IVSVTX4 U484 ( .A(num_i[11]), .Z(n190) );
  ND2SVTX8 U485 ( .A(n478), .B(n469), .Z(n442) );
  NR2SVTX8 U486 ( .A(num_i[24]), .B(num_i[25]), .Z(n469) );
  NR2SVTX8 U487 ( .A(num_i[27]), .B(num_i[26]), .Z(n478) );
  IVSVTX12 U488 ( .A(n442), .Z(n399) );
  IVSVTX4 U489 ( .A(n195), .Z(n372) );
  ND4SVTX4 U490 ( .A(n353), .B(n493), .C(n195), .D(n289), .Z(n288) );
  ND4ABSVTX8 U491 ( .A(n489), .B(n490), .C(n287), .D(n286), .Z(n195) );
  CTIVSVTX4 U492 ( .A(n198), .Z(n407) );
  AO7ABSVTX8 U493 ( .A(n587), .B(n570), .C(n228), .Z(n571) );
  IVSVTX10 U494 ( .A(n727), .Z(n246) );
  IVSVTX4 U495 ( .A(rslt_o[31]), .Z(n196) );
  ND3SVTX6 U496 ( .A(n196), .B(n657), .C(n586), .Z(n350) );
  ND2SVTX4 U497 ( .A(n711), .B(n217), .Z(n637) );
  IVSVTX4 U498 ( .A(n600), .Z(n602) );
  BFSVTX12 U499 ( .A(n419), .Z(n309) );
  AO2SVTX6 U500 ( .A(n292), .B(num_i[11]), .C(n301), .D(n603), .Z(n543) );
  IVSVTX10 U501 ( .A(n679), .Z(n271) );
  BFSVTX2 U502 ( .A(n449), .Z(n226) );
  IVSVTX4 U503 ( .A(n703), .Z(n197) );
  AO2SVTX8 U504 ( .A(n548), .B(n327), .C(n567), .D(n471), .Z(n651) );
  IVSVTX8 U505 ( .A(n306), .Z(n304) );
  AO4SVTX4 U506 ( .A(n346), .B(n333), .C(n713), .D(n199), .Z(n223) );
  NR2SVTX4 U507 ( .A(n367), .B(n536), .Z(n341) );
  ND2SVTX4 U508 ( .A(n228), .B(n453), .Z(n198) );
  ND2SVTX4 U509 ( .A(n684), .B(n200), .Z(n546) );
  NR2SVTX4 U510 ( .A(n187), .B(n594), .Z(n200) );
  ND3ASVTX6 U511 ( .A(n693), .B(n362), .C(n361), .Z(n256) );
  IVSVTX4 U512 ( .A(num_i[21]), .Z(n517) );
  ND3ABSVTX8 U513 ( .A(num_i[21]), .B(num_i[20]), .C(n231), .Z(n413) );
  CTIVSVTX8 U514 ( .A(n409), .Z(n477) );
  ND2SVTX6 U515 ( .A(n362), .B(n361), .Z(n217) );
  AO7SVTX4 U516 ( .A(n301), .B(n646), .C(n645), .Z(n649) );
  AO7SVTX8 U517 ( .A(n679), .B(n462), .C(n398), .Z(n440) );
  AO7ABSVTX8 U518 ( .A(n202), .B(n718), .C(n294), .Z(n636) );
  NR2ASVTX6 U519 ( .A(n706), .B(rslt_o[31]), .Z(n202) );
  IVSVTX8 U520 ( .A(n218), .Z(n227) );
  ND2SVTX6 U521 ( .A(n277), .B(n665), .Z(n414) );
  ND2SVTX4 U522 ( .A(n695), .B(n694), .Z(n696) );
  AO1SVTX8 U523 ( .A(n246), .B(n642), .C(n214), .D(n269), .Z(n203) );
  ND2ASVTX8 U524 ( .A(n303), .B(n449), .Z(n411) );
  ND2ASVTX8 U525 ( .A(n204), .B(n399), .Z(n449) );
  IVSVTX4 U526 ( .A(n413), .Z(n204) );
  IVSVTX4 U527 ( .A(n589), .Z(n343) );
  ND2ASVTX8 U528 ( .A(n644), .B(n643), .Z(keyvalues_m1[18]) );
  AO2SVTX6 U529 ( .A(n273), .B(n599), .C(n396), .D(n684), .Z(n205) );
  ND2SVTX4 U530 ( .A(num_i[3]), .B(n471), .Z(n552) );
  IVSVTX4 U531 ( .A(n206), .Z(n548) );
  ND2SVTX4 U532 ( .A(num_i[10]), .B(n227), .Z(n206) );
  BFSVTX1 U533 ( .A(n544), .Z(n207) );
  ND2SVTX4 U534 ( .A(n438), .B(n383), .Z(n362) );
  IVSVTX4 U535 ( .A(n694), .Z(n312) );
  IVSVTX8 U536 ( .A(n230), .Z(n446) );
  AO7SVTX6 U537 ( .A(n207), .B(n718), .C(n545), .Z(n684) );
  AO7SVTX6 U538 ( .A(n711), .B(n726), .C(n209), .Z(n208) );
  IVSVTX4 U539 ( .A(n414), .Z(n451) );
  AO4SVTX4 U540 ( .A(n210), .B(n271), .C(n702), .D(n727), .Z(keyvalues_m1[9])
         );
  ND3SVTX8 U541 ( .A(n575), .B(n320), .C(n189), .Z(n318) );
  ND4SVTX6 U542 ( .A(n492), .B(n371), .C(n368), .D(n370), .Z(n353) );
  NR2SVTX6 U543 ( .A(num_i[31]), .B(num_i[30]), .Z(n406) );
  AO7ABSVTX8 U544 ( .A(n336), .B(n699), .C(n701), .Z(n335) );
  AO4SVTX4 U545 ( .A(n594), .B(n690), .C(n661), .D(n279), .Z(n211) );
  NR2SVTX4 U546 ( .A(n620), .B(n228), .Z(n431) );
  IVSVTX12 U547 ( .A(n467), .Z(n703) );
  IVSVTX6 U548 ( .A(n467), .Z(n218) );
  MUX21NSVTX6 U549 ( .A(n642), .B(n284), .S(n711), .Z(n643) );
  AO6SVTX4 U550 ( .A(n453), .B(n691), .C(n590), .Z(n593) );
  NR2SVTX4 U551 ( .A(n710), .B(n727), .Z(n425) );
  ND2SVTX4 U552 ( .A(n721), .B(n213), .Z(n212) );
  AO6SVTX8 U553 ( .A(n385), .B(n712), .C(n268), .Z(n214) );
  NR2SVTX8 U554 ( .A(n380), .B(n372), .Z(n355) );
  ND2SVTX6 U555 ( .A(n651), .B(n305), .Z(n549) );
  IVSVTX4 U556 ( .A(n215), .Z(n269) );
  ND2ASVTX8 U557 ( .A(n249), .B(n462), .Z(n432) );
  AO7SVTX4 U558 ( .A(n454), .B(n713), .C(n641), .Z(n644) );
  AO6SVTX8 U559 ( .A(n256), .B(n255), .C(n253), .Z(n444) );
  AO7SVTX2 U560 ( .A(n709), .B(n534), .C(n630), .Z(n631) );
  AO6SVTX6 U561 ( .A(n575), .B(num_i[14]), .C(n455), .Z(n528) );
  NR3SVTX8 U562 ( .A(n463), .B(n584), .C(n663), .Z(n677) );
  IVSVTX4 U563 ( .A(n681), .Z(n682) );
  ND2SVTX4 U564 ( .A(n635), .B(n416), .Z(n547) );
  F_MUX21SVTX6 U565 ( .A(n576), .B(n706), .S(n693), .Z(n565) );
  ND3SVTX8 U566 ( .A(n434), .B(n228), .C(n306), .Z(n694) );
  NR2SVTX4 U567 ( .A(n535), .B(n340), .Z(n700) );
  ND2SVTX4 U568 ( .A(n633), .B(n383), .Z(n221) );
  IVSVTX8 U569 ( .A(n222), .Z(n453) );
  NR2SVTX4 U570 ( .A(n532), .B(n531), .Z(n222) );
  ND3ASVTX8 U571 ( .A(n457), .B(n527), .C(n353), .Z(n380) );
  ND3ABSVTX6 U572 ( .A(n228), .B(n283), .C(n364), .Z(n262) );
  AO6SVTX8 U573 ( .A(rslt_o[31]), .B(n569), .C(n568), .Z(n283) );
  OR2SVTX8 U574 ( .A(n297), .B(n442), .Z(n467) );
  IVSVTX4 U575 ( .A(n354), .Z(n275) );
  ND2ASVTX8 U576 ( .A(n676), .B(n364), .Z(n720) );
  ND2SVTX4 U577 ( .A(n438), .B(n347), .Z(n556) );
  AO3SVTX4 U578 ( .A(n604), .B(n529), .C(n616), .D(n491), .Z(n527) );
  IVSVTX10 U579 ( .A(n354), .Z(n279) );
  ND3SVTX6 U580 ( .A(n249), .B(n678), .C(n298), .Z(n680) );
  IVSVTX8 U581 ( .A(n227), .Z(n463) );
  ND3SVTX6 U582 ( .A(n647), .B(n703), .C(n183), .Z(n587) );
  ND2SVTX8 U583 ( .A(n252), .B(n251), .Z(n306) );
  AO7SVTX8 U584 ( .A(n588), .B(n446), .C(n587), .Z(n434) );
  ND2SVTX4 U585 ( .A(n693), .B(n402), .Z(n315) );
  AO7SVTX6 U586 ( .A(n451), .B(n696), .C(n693), .Z(n697) );
  AO2SVTX8 U587 ( .A(n314), .B(n670), .C(n313), .D(n225), .Z(keyvalues_m1[14])
         );
  IVSVTX12 U588 ( .A(n234), .Z(keyvalues_m1[27]) );
  ND2ASVTX8 U589 ( .A(n237), .B(n235), .Z(n234) );
  NR2SVTX4 U590 ( .A(rslt_o[27]), .B(n239), .Z(n237) );
  AO2SVTX6 U591 ( .A(n179), .B(n328), .C(n238), .D(n246), .Z(keyvalues_m1[26])
         );
  ND2SVTX4 U592 ( .A(n388), .B(n478), .Z(n325) );
  IVSVTX12 U593 ( .A(n240), .Z(n693) );
  NR3ABSVTX8 U594 ( .A(n241), .B(n177), .C(n408), .Z(n240) );
  ND3SVTX8 U595 ( .A(n243), .B(n242), .C(n244), .Z(n408) );
  ND3SVTX8 U596 ( .A(n502), .B(n503), .C(n188), .Z(n242) );
  IVSVTX4 U597 ( .A(n727), .Z(n711) );
  BFSVTX6 U598 ( .A(n408), .Z(n249) );
  ND2SVTX4 U599 ( .A(n481), .B(n191), .Z(n516) );
  ND3SVTX8 U600 ( .A(n376), .B(n355), .C(n374), .Z(n531) );
  AO7ABSVTX4 U601 ( .A(n416), .B(n714), .C(n254), .Z(n253) );
  ND2SVTX4 U602 ( .A(n396), .B(n715), .Z(n254) );
  OR3ABCSVTX6 U603 ( .A(n578), .B(n703), .C(n183), .Z(n600) );
  ND3SVTX8 U604 ( .A(n540), .B(n357), .C(n356), .Z(n609) );
  IVSVTX4 U605 ( .A(n306), .Z(n367) );
  ND3SVTX8 U606 ( .A(n342), .B(n262), .C(n270), .Z(n642) );
  ND4SVTX4 U607 ( .A(num_i[25]), .B(n492), .C(n616), .D(n194), .Z(n495) );
  IVSVTX4 U608 ( .A(n266), .Z(n545) );
  IVSVTX8 U609 ( .A(n727), .Z(n268) );
  NR2SVTX6 U610 ( .A(num_i[29]), .B(num_i[28]), .Z(n370) );
  ND2ASVTX8 U611 ( .A(n257), .B(n275), .Z(n274) );
  IVSVTX8 U612 ( .A(n181), .Z(n276) );
  AO6ASVTX8 U613 ( .A(n663), .B(n435), .C(n280), .Z(n653) );
  IVSVTX4 U614 ( .A(n551), .Z(n280) );
  AO7SVTX8 U615 ( .A(n476), .B(n283), .C(n664), .Z(n665) );
  ND2SVTX6 U616 ( .A(n388), .B(n387), .Z(n523) );
  NR2SVTX4 U617 ( .A(n523), .B(n442), .Z(n378) );
  ND2SVTX4 U618 ( .A(n624), .B(n345), .Z(n623) );
  IVSVTX4 U619 ( .A(rslt_o[31]), .Z(n624) );
  NR3SVTX8 U620 ( .A(n520), .B(n488), .C(n330), .Z(n286) );
  NR3SVTX8 U621 ( .A(n487), .B(n455), .C(n486), .Z(n287) );
  ND3SVTX8 U622 ( .A(n189), .B(n291), .C(n418), .Z(n497) );
  NR2SVTX8 U623 ( .A(n538), .B(n334), .Z(n418) );
  IVSVTX6 U624 ( .A(num_i[20]), .Z(n295) );
  ND2SVTX8 U625 ( .A(n510), .B(n663), .Z(n718) );
  ND2SVTX8 U626 ( .A(n296), .B(n496), .Z(n303) );
  NR2SVTX8 U627 ( .A(num_i[31]), .B(num_i[30]), .Z(n496) );
  NR2SVTX6 U628 ( .A(num_i[28]), .B(num_i[29]), .Z(n296) );
  ND3ABSVTX6 U629 ( .A(num_i[28]), .B(num_i[29]), .C(n496), .Z(n297) );
  ND3SVTX6 U630 ( .A(n272), .B(n678), .C(n298), .Z(n553) );
  AO6CSVTX8 U631 ( .A(n347), .B(n685), .C(n405), .Z(n299) );
  NR2SVTX6 U632 ( .A(n532), .B(n531), .Z(n300) );
  ND2SVTX4 U633 ( .A(n617), .B(n467), .Z(n645) );
  IVSVTX8 U634 ( .A(num_i[28]), .Z(n616) );
  IVSVTX8 U635 ( .A(num_i[29]), .Z(n491) );
  ND2SVTX4 U636 ( .A(n365), .B(n308), .Z(n307) );
  IVSVTX12 U637 ( .A(n693), .Z(n727) );
  ND2SVTX6 U638 ( .A(n187), .B(n316), .Z(n402) );
  NR2SVTX8 U639 ( .A(n692), .B(n279), .Z(n316) );
  ND3SVTX8 U640 ( .A(n228), .B(n366), .C(n277), .Z(n317) );
  ND2SVTX6 U641 ( .A(n697), .B(n381), .Z(keyvalues_m1[13]) );
  NR2SVTX2 U642 ( .A(num_i[28]), .B(num_i[29]), .Z(n332) );
  ND2SVTX8 U643 ( .A(n323), .B(n322), .Z(n331) );
  NR2SVTX6 U644 ( .A(num_i[28]), .B(num_i[30]), .Z(n322) );
  NR2SVTX8 U645 ( .A(num_i[31]), .B(num_i[29]), .Z(n323) );
  ND2SVTX4 U646 ( .A(n387), .B(n469), .Z(n324) );
  ND2ASVTX8 U647 ( .A(n331), .B(n418), .Z(n522) );
  IVSVTX4 U648 ( .A(n539), .Z(n326) );
  MUX21NSVTX6 U649 ( .A(n677), .B(n676), .S(n279), .Z(n717) );
  AO7ABSVTX4 U650 ( .A(n416), .B(n438), .C(n329), .Z(n683) );
  NR2SVTX4 U651 ( .A(n373), .B(n331), .Z(n379) );
  ND2SVTX4 U652 ( .A(n404), .B(n279), .Z(n403) );
  ND2SVTX6 U653 ( .A(n703), .B(n183), .Z(n559) );
  ND2SVTX4 U654 ( .A(n640), .B(n271), .Z(n333) );
  AO4SVTX6 U655 ( .A(n559), .B(n481), .C(n463), .D(n207), .Z(n640) );
  ND4ABSVTX8 U656 ( .A(n506), .B(n334), .C(n505), .D(n412), .Z(n540) );
  ND2SVTX6 U657 ( .A(n478), .B(n469), .Z(n334) );
  ND2SVTX8 U658 ( .A(n338), .B(n339), .Z(keyvalues_m1[23]) );
  NR2ASVTX6 U659 ( .A(num_i[11]), .B(n703), .Z(n655) );
  NR2SVTX8 U660 ( .A(n532), .B(n531), .Z(n354) );
  ND2SVTX4 U661 ( .A(n434), .B(n343), .Z(n342) );
  AO17SVTX4 U662 ( .A(n608), .B(n345), .C(n607), .D(n228), .Z(n613) );
  NR2SVTX2 U663 ( .A(n523), .B(n539), .Z(n509) );
  NR3ABSVTX8 U664 ( .A(n192), .B(n190), .C(n516), .Z(n539) );
  ND2ASVTX8 U665 ( .A(n464), .B(n594), .Z(n346) );
  ND2SVTX4 U666 ( .A(n348), .B(n383), .Z(n360) );
  NR2SVTX6 U667 ( .A(num_i[24]), .B(num_i[25]), .Z(n485) );
  ND3SVTX6 U668 ( .A(rslt_o[29]), .B(n555), .C(n364), .Z(n533) );
  ND2SVTX4 U669 ( .A(n662), .B(n365), .Z(n650) );
  ND2SVTX4 U670 ( .A(n591), .B(n304), .Z(n592) );
  NR2SVTX4 U671 ( .A(num_i[25]), .B(n369), .Z(n368) );
  IVSVTX4 U672 ( .A(num_i[23]), .Z(n369) );
  NR2SVTX4 U673 ( .A(num_i[24]), .B(num_i[30]), .Z(n371) );
  ND2SVTX6 U674 ( .A(n477), .B(n375), .Z(n374) );
  ND2SVTX4 U675 ( .A(n417), .B(n382), .Z(n381) );
  ND3SVTX8 U676 ( .A(n563), .B(n564), .C(n562), .Z(keyvalues_m1[21]) );
  ND2ASVTX8 U677 ( .A(n384), .B(n273), .Z(n671) );
  NR2SVTX4 U678 ( .A(n591), .B(n228), .Z(n404) );
  NR3SVTX8 U679 ( .A(n687), .B(n386), .C(n428), .Z(n674) );
  AO6CSVTX6 U680 ( .A(n473), .B(n419), .C(n194), .Z(n626) );
  ND2SVTX4 U681 ( .A(n272), .B(n702), .Z(n398) );
  ND2SVTX6 U682 ( .A(n705), .B(n565), .Z(n566) );
  MUX21NSVTX8 U683 ( .A(n410), .B(n704), .S(n305), .Z(n722) );
  NR3SVTX6 U684 ( .A(n728), .B(n463), .C(n464), .Z(n410) );
  NR2SVTX4 U685 ( .A(n228), .B(n305), .Z(n415) );
  AO17SVTX8 U686 ( .A(n574), .B(n425), .C(n424), .D(n582), .Z(keyvalues_m1[15]) );
  NR2ASVTX6 U687 ( .A(n426), .B(n631), .Z(n632) );
  ND2SVTX6 U688 ( .A(n638), .B(n637), .Z(keyvalues_m1[19]) );
  ND2SVTX4 U689 ( .A(n464), .B(n438), .Z(n536) );
  ND2SVTX4 U690 ( .A(rslt_o[28]), .B(n427), .Z(n699) );
  AO7ABSVTX8 U691 ( .A(n542), .B(n347), .C(n541), .Z(n428) );
  ND3SVTX6 U692 ( .A(n430), .B(n429), .C(n178), .Z(n634) );
  IVSVTX4 U693 ( .A(n621), .Z(n429) );
  NR2SVTX4 U694 ( .A(n622), .B(n431), .Z(n430) );
  ND2SVTX4 U695 ( .A(n517), .B(n295), .Z(n488) );
  IVSVTX12 U696 ( .A(n433), .Z(keyvalues_m1[12]) );
  ND2SVTX4 U697 ( .A(n653), .B(n453), .Z(n678) );
  AO2SVTX6 U698 ( .A(n292), .B(n625), .C(n301), .D(n520), .Z(n437) );
  IVSVTX12 U699 ( .A(n440), .Z(keyvalues_m1[10]) );
  ND2SVTX4 U700 ( .A(n687), .B(n441), .Z(n562) );
  ND2SVTX4 U701 ( .A(n466), .B(n700), .Z(n701) );
  IVSVTX12 U702 ( .A(n443), .Z(keyvalues_m1[8]) );
  IVSVTX12 U703 ( .A(n444), .Z(n445) );
  AO7SVTX6 U704 ( .A(n452), .B(n722), .C(n708), .Z(keyvalues_m1[2]) );
  MUX21NSVTX8 U705 ( .A(n716), .B(n723), .S(n272), .Z(keyvalues_m1[4]) );
  ND2SVTX2 U706 ( .A(n579), .B(n183), .Z(n580) );
  OR2SVTX4 U707 ( .A(n539), .B(n538), .Z(n447) );
  NR2SVTX4 U708 ( .A(num_i[16]), .B(num_i[17]), .Z(n482) );
  ND3ASVTX2 U709 ( .A(n191), .B(n327), .C(n301), .Z(n550) );
  IVSVTX12 U710 ( .A(n460), .Z(keyvalues_m1[16]) );
  BFSVTX4 U711 ( .A(num_i[29]), .Z(n526) );
  MUX21NSVTX8 U712 ( .A(n583), .B(n704), .S(n594), .Z(n716) );
  AO21SVTX8 U713 ( .A(n679), .B(n719), .C(n554), .D(n553), .Z(keyvalues_m1[7])
         );
  AO7SVTX8 U714 ( .A(n673), .B(n672), .C(n246), .Z(n564) );
  BFSVTX10 U715 ( .A(num_i[22]), .Z(n520) );
  IVSVTX4 U716 ( .A(n504), .Z(n465) );
  ND2ASVTX1 U717 ( .A(n707), .B(n679), .Z(n708) );
  ND3SVTX4 U718 ( .A(n272), .B(n549), .C(n720), .Z(n721) );
  ND2ASVTX1 U719 ( .A(n464), .B(n594), .Z(n454) );
  MUX21NSVTX8 U720 ( .A(n716), .B(n717), .S(n249), .Z(keyvalues_m1[5]) );
  AO6CSVTX4 U721 ( .A(n194), .B(n526), .C(n456), .Z(n493) );
  IVSVTX12 U722 ( .A(n453), .Z(n594) );
  ND3SVTX1 U723 ( .A(n399), .B(n576), .C(n506), .Z(n577) );
  ND3ABSVTX4 U724 ( .A(n710), .B(n271), .C(n574), .Z(n459) );
  ND2SVTX4 U725 ( .A(n396), .B(n714), .Z(n641) );
  OR2SVTX4 U726 ( .A(n186), .B(n713), .Z(n475) );
  AO7SVTX2 U727 ( .A(n192), .B(rslt_o[31]), .C(n530), .Z(n633) );
  ND2ASVTX1 U728 ( .A(n192), .B(n471), .Z(n664) );
  ND3SVTX4 U729 ( .A(n604), .B(n616), .C(n194), .Z(n494) );
  BFSVTX2 U730 ( .A(num_i[15]), .Z(n578) );
  NR3SVTX6 U731 ( .A(n646), .B(n463), .C(n464), .Z(n585) );
  ND2SVTX4 U732 ( .A(n396), .B(n636), .Z(n557) );
  IVSVTX2 U733 ( .A(n511), .Z(n512) );
  NR2SVTX2 U734 ( .A(n455), .B(n544), .Z(n484) );
  AN2SVTX8 U735 ( .A(n580), .B(n581), .Z(n691) );
  AO7SVTX4 U736 ( .A(rslt_o[31]), .B(n191), .C(n620), .Z(n555) );
  IVSVTX8 U737 ( .A(n184), .Z(n618) );
  ND2SVTX4 U738 ( .A(n578), .B(n227), .Z(n581) );
  NR2ASVTX4 U739 ( .A(n576), .B(n183), .Z(n608) );
  ND2SVTX4 U740 ( .A(n725), .B(n724), .Z(n726) );
  NR2SVTX2 U741 ( .A(num_i[25]), .B(num_i[27]), .Z(n521) );
  ND2SVTX4 U742 ( .A(n181), .B(n273), .Z(n582) );
  ND2SVTX2 U743 ( .A(n596), .B(n227), .Z(n537) );
  AN2SVTX8 U744 ( .A(n508), .B(n309), .Z(n471) );
  AN2SVTX4 U745 ( .A(n663), .B(n226), .Z(n476) );
  AN3CSVTX8 U746 ( .A(n703), .B(num_i[3]), .C(n477), .Z(n654) );
  BFSVTX12 U747 ( .A(n183), .Z(rslt_o[31]) );
  AN3SVTX1 U748 ( .A(n506), .B(n399), .C(n657), .Z(n472) );
  IVSVTX4 U749 ( .A(n665), .Z(n668) );
  BFSVTX2 U750 ( .A(num_i[14]), .Z(n625) );
  NR2SVTX6 U751 ( .A(num_i[19]), .B(num_i[17]), .Z(n479) );
  ND3ABSVTX8 U752 ( .A(num_i[16]), .B(num_i[18]), .C(n479), .Z(n506) );
  BFSVTX2 U753 ( .A(num_i[21]), .Z(n596) );
  AO17SVTX4 U754 ( .A(n501), .B(n728), .C(n500), .D(n499), .Z(n503) );
  AO6SVTX4 U755 ( .A(n188), .B(n509), .C(n508), .Z(n510) );
  NR2SVTX2 U756 ( .A(num_i[2]), .B(num_i[3]), .Z(n511) );
  ND2SVTX4 U757 ( .A(n513), .B(n512), .Z(n515) );
  AO6CSVTX2 U758 ( .A(n703), .B(n487), .C(n519), .Z(n620) );
  BFSVTX1 U759 ( .A(num_i[23]), .Z(n601) );
  ND3SVTX2 U760 ( .A(n369), .B(n600), .C(n561), .Z(n542) );
  AO7ABSVTX4 U761 ( .A(n706), .B(n471), .C(n550), .Z(n676) );
  NR2ASVTX6 U762 ( .A(n567), .B(n301), .Z(n569) );
  ND2SVTX4 U763 ( .A(n667), .B(n464), .Z(n572) );
  ND2SVTX4 U764 ( .A(n487), .B(n618), .Z(n570) );
  ND2SVTX6 U765 ( .A(n572), .B(n571), .Z(n573) );
  NR2SVTX4 U766 ( .A(n658), .B(n472), .Z(n591) );
  AO7SVTX2 U767 ( .A(n185), .B(rslt_o[31]), .C(n450), .Z(n595) );
  IVSVTX0H U768 ( .A(n603), .Z(n606) );
  IVSVTX0H U769 ( .A(n604), .Z(n605) );
  AO7SVTX2 U770 ( .A(n301), .B(n295), .C(n616), .Z(n622) );
  F_ND2ASVTX2 U771 ( .A(n349), .B(n471), .Z(n652) );
  ND2SVTX4 U772 ( .A(n662), .B(n277), .Z(n725) );
  ND2ASVTX8 U773 ( .A(n367), .B(n668), .Z(n724) );
  NR3SVTX8 U774 ( .A(n673), .B(rslt_o[27]), .C(n672), .Z(n675) );
  AO7SVTX8 U775 ( .A(n674), .B(n675), .C(n475), .Z(keyvalues_m1[22]) );
  NR2SVTX4 U776 ( .A(n698), .B(n686), .Z(n688) );
endmodule

